`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:50:28 01/03/2019 
// Design Name: 
// Module Name:    pipesmod 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pipesmod(input wire [9:0] x,
                input wire [9:0] y,
                input wire [3:0]mode,  // 0-7 are pipes, 8 and 9 are the starting and ending points pixel val
					 output wire [11:0]out
                );	 
	reg [11:0]data[0:63999] = {
// pipe zero horizontal straight pipe

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hccc, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hbbb, 12'hccc, 12'hbbb, 12'hccc, 12'hddd, 12'hfff, 12'h777, 
12'h888, 12'h888, 12'h666, 12'h888, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'h999, 12'h777, 12'h777, 12'h888, 12'h888, 12'h666, 12'h888, 12'hddd, 12'h333, 
12'h444, 12'h444, 12'h222, 12'h222, 12'h777, 12'haaa, 12'haaa, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h777, 12'h444, 12'h333, 12'h444, 12'h444, 12'h000, 12'h333, 12'hbbb, 12'h888, 
12'h888, 12'h999, 12'h888, 12'h555, 12'h555, 12'haaa, 12'hbbb, 12'haaa, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h666, 12'h555, 12'hbbb, 12'heee, 
12'heee, 12'heee, 12'hddd, 12'h888, 12'h777, 12'hddd, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'haaa, 12'haaa, 12'hddd, 12'heee, 12'haaa, 12'h888, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'h777, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'h999, 12'h777, 12'hbbb, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hccc, 12'h999, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'h999, 12'h555, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'h777, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'h999, 12'h333, 12'h777, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h222, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'h999, 12'h666, 12'h777, 12'h777, 12'h555, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h555, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h555, 12'h666, 12'h888, 12'h444, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h999, 12'hccc, 12'hccc, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hddd, 12'h888, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h888, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'h777, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hbbb, 12'hddd, 
12'hddd, 12'hddd, 12'hccc, 12'h888, 12'h555, 12'h888, 12'haaa, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'haaa, 12'h555, 12'h666, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h777, 12'hbbb, 12'h777, 
12'h777, 12'h777, 12'h666, 12'h444, 12'h777, 12'hbbb, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'haaa, 12'hccc, 12'hccc, 12'h888, 12'h444, 12'h666, 12'h777, 12'h777, 12'h777, 12'h555, 12'h555, 12'hbbb, 12'h111, 
12'h000, 12'h000, 12'h111, 12'h000, 12'h888, 12'hddd, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'h000, 
12'h111, 12'h111, 12'h111, 12'h222, 12'h666, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'h777, 12'h444, 12'h222, 12'h111, 12'h111, 12'h111, 12'h000, 12'h555, 12'hccc, 12'h000, 
12'h111, 12'h000, 12'h222, 12'h333, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h333, 12'h333, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h555, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h333, 12'h444, 12'h444, 12'h333, 12'h222, 12'h333, 12'h444, 12'h444, 12'h333, 12'h111, 12'h111, 12'h111, 12'h000, 12'h555, 12'hccc, 12'h000, 
12'h000, 12'h000, 12'h000, 12'h333, 12'h222, 12'h111, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h555, 12'hccc, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h555, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h222, 12'h333, 12'h333, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h444, 12'h555, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'hccc, 12'haaa, 
12'hbbb, 12'hbbb, 12'haaa, 12'h777, 12'h444, 12'h555, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h333, 12'h666, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'h666, 12'hbbb, 12'hddd, 
12'hddd, 12'hddd, 12'hccc, 12'h888, 12'h666, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h666, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h777, 12'hbbb, 12'hccc, 
12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h666, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'hbbb, 12'hccc, 
12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h666, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'hbbb, 12'hccc, 
12'hccc, 12'hddd, 12'hccc, 12'h888, 12'h666, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'hbbb, 12'hccc, 
12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h666, 12'h888, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h555, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'hbbb, 12'hccc, 
12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h555, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'h444, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'hbbb, 12'hccc, 
12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h666, 12'hbbb, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'haaa, 12'hbbb, 12'hccc, 12'h777, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'hbbb, 12'hccc, 
12'hccc, 12'hccc, 12'hbbb, 12'h666, 12'h777, 12'hddd, 12'heee, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hddd, 12'heee, 12'h888, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'hbbb, 12'haaa, 
12'hbbb, 12'hbbb, 12'haaa, 12'h666, 12'h777, 12'hbbb, 12'hccc, 12'haaa, 12'h888, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'h777, 12'h555, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'h666, 12'hbbb, 12'h999, 
12'haaa, 12'h999, 12'h999, 12'h666, 12'h555, 12'h777, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h777, 12'h555, 12'h555, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h777, 12'h666, 12'hbbb, 12'haaa, 
12'haaa, 12'haaa, 12'h999, 12'h666, 12'h444, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h444, 12'h555, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h666, 12'hbbb, 12'haaa, 
12'haaa, 12'haaa, 12'h999, 12'h777, 12'h666, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h666, 12'h666, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h666, 12'hbbb, 12'haaa, 
12'haaa, 12'haaa, 12'h999, 12'h666, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'h666, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h666, 12'hbbb, 12'h999, 
12'haaa, 12'haaa, 12'h999, 12'h666, 12'h888, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'h888, 12'h666, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h666, 12'hbbb, 12'h999, 
12'haaa, 12'haaa, 12'h999, 12'h666, 12'h777, 12'haaa, 12'hbbb, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'hbbb, 12'h888, 12'h555, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h666, 12'hbbb, 12'hbbb, 
12'hbbb, 12'hbbb, 12'haaa, 12'h666, 12'h777, 12'hccc, 12'hddd, 12'hbbb, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'hbbb, 12'haaa, 12'hccc, 12'hddd, 12'h777, 12'h555, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'h888, 12'h666, 12'hbbb, 12'heee, 
12'heee, 12'heee, 12'hddd, 12'h777, 12'h666, 12'hccc, 12'heee, 12'hbbb, 12'h888, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h888, 12'haaa, 12'hddd, 12'hddd, 12'h777, 12'h666, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'h777, 12'hbbb, 12'heee, 
12'heee, 12'hfff, 12'hddd, 12'h777, 12'h777, 12'hccc, 12'hddd, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hddd, 12'h777, 12'h555, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h666, 12'haaa, 12'heee, 
12'heee, 12'heee, 12'hddd, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h888, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h888, 12'hccc, 12'heee, 
12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'heee, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 

// pipe one, vertical straight pipe



12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h888, 12'h888, 12'h888, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h888, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h444, 12'h000, 12'h111, 12'h111, 12'h000, 12'h666, 12'haaa, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hbbb, 12'h666, 12'h000, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'haaa, 12'h666, 12'h000, 12'h000, 12'h000, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h333, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h666, 12'h000, 12'h111, 12'h111, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h666, 12'h000, 12'h111, 12'h111, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hccc, 12'haaa, 12'h666, 12'h000, 12'h222, 12'h111, 12'h000, 12'h777, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'h888, 12'h222, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h555, 12'h333, 12'h333, 12'h222, 12'h000, 12'h444, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h888, 12'h555, 12'h333, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'h666, 12'h777, 12'h777, 12'h888, 12'h777, 12'h666, 12'h444, 12'h555, 12'h777, 12'h777, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h444, 12'h222, 12'h222, 12'h333, 12'h666, 12'h888, 12'h777, 12'h555, 12'h888, 12'h999, 12'h666, 12'h333, 12'h555, 12'h777, 12'h777, 12'h555, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'hbbb, 12'hbbb, 12'h999, 12'h777, 12'h777, 12'hbbb, 12'hddd, 12'hbbb, 12'h777, 12'h888, 12'h999, 12'h888, 12'h888, 12'h999, 12'h555, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hbbb, 12'h888, 12'haaa, 12'hccc, 12'h777, 12'h777, 12'haaa, 12'hbbb, 12'hddd, 12'haaa, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'heee, 12'hddd, 12'hbbb, 12'hddd, 12'heee, 12'hccc, 12'hbbb, 12'h999, 12'hccc, 12'heee, 12'hccc, 12'h888, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'h777, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hccc, 12'haaa, 12'hddd, 12'hccc, 12'h777, 12'haaa, 12'hddd, 12'hccc, 12'heee, 12'hbbb, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'heee, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h333, 12'h999, 12'hbbb, 12'haaa, 12'hbbb, 12'heee, 12'haaa, 12'h555, 12'haaa, 12'heee, 12'hbbb, 12'hbbb, 12'haaa, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'haaa, 12'heee, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h111, 12'h000, 12'h333, 12'haaa, 12'h999, 12'haaa, 12'heee, 12'hfff, 12'hbbb, 12'h444, 12'haaa, 12'hfff, 12'hddd, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h444, 12'hccc, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h333, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h333, 12'h111, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h222, 12'h111, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h111, 12'h000, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h333, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'hbbb, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'hbbb, 12'heee, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h111, 12'h000, 12'h444, 12'hbbb, 12'h999, 12'hbbb, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'heee, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h111, 12'h000, 12'h333, 12'h999, 12'hbbb, 12'haaa, 12'hccc, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'heee, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hddd, 12'hccc, 12'haaa, 12'hddd, 12'hfff, 12'hddd, 12'hbbb, 12'h999, 12'hbbb, 12'hddd, 12'hbbb, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h333, 12'h999, 12'hddd, 12'hccc, 12'haaa, 12'hddd, 12'hbbb, 12'h666, 12'haaa, 12'hddd, 12'hbbb, 12'hddd, 12'haaa, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'hccc, 12'hccc, 12'haaa, 12'h888, 12'h777, 12'hccc, 12'heee, 12'hccc, 12'h777, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h666, 12'h111, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hccc, 12'haaa, 12'hccc, 12'hddd, 12'h888, 12'h888, 12'hccc, 12'hccc, 12'heee, 12'haaa, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h666, 12'h444, 12'h555, 12'h777, 12'h888, 12'h777, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h333, 12'h333, 12'h333, 12'h444, 12'h777, 12'h999, 12'h888, 12'h555, 12'h777, 12'h888, 12'h444, 12'h222, 12'h777, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h555, 12'h666, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h444, 12'h444, 12'h444, 12'h444, 12'h333, 12'h444, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h999, 12'h888, 12'h888, 12'h777, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'h999, 12'h555, 12'h000, 12'h222, 12'h222, 12'h000, 12'h666, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h888, 12'h444, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h666, 12'h111, 12'h111, 12'h000, 12'h111, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h333, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h666, 12'h000, 12'h111, 12'h111, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h666, 12'h000, 12'h111, 12'h111, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'h999, 12'h555, 12'h000, 12'h000, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h666, 12'h111, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 



// pipe two, left to bottom 90 degrees

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 
12'hccc, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h666, 12'h666, 12'h777, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 
12'h222, 12'h444, 12'h333, 12'h666, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 
12'h777, 12'h888, 12'h555, 12'h777, 12'hbbb, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hddd, 12'heee, 12'haaa, 12'h999, 12'hccc, 12'hbbb, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hfff, 12'hfff, 12'hccc, 12'h888, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'hccc, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'hccc, 12'h666, 12'h999, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'hccc, 12'h777, 12'h555, 12'h444, 12'h444, 12'h444, 12'h555, 12'h666, 12'h777, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'hccc, 12'haaa, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h666, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hfff, 12'hfff, 12'hccc, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h555, 12'h444, 12'h444, 12'h666, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hddd, 12'heee, 12'hbbb, 12'h666, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'haaa, 12'h888, 12'h666, 12'h444, 12'h555, 12'h777, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 
12'h555, 12'h666, 12'h333, 12'h888, 12'hccc, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h666, 12'h444, 12'h444, 12'h666, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 
12'h111, 12'h000, 12'h000, 12'h999, 12'hddd, 12'hbbb, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h777, 12'h555, 12'h444, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 
12'h000, 12'h000, 12'h111, 12'h777, 12'haaa, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h444, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 
12'h111, 12'h111, 12'h333, 12'h444, 12'h444, 12'h555, 12'h888, 12'h888, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h333, 12'h555, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 
12'h111, 12'h111, 12'h333, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h666, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h555, 12'h222, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 
12'h444, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'h333, 12'h666, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h888, 12'h555, 12'h666, 12'h666, 12'h555, 12'h444, 12'h444, 12'h444, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h222, 12'h555, 12'h999, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h444, 12'h444, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hccc, 12'hddd, 12'haaa, 12'h777, 12'haaa, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h777, 12'h555, 12'h333, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h555, 12'h444, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hddd, 12'haaa, 12'h777, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h555, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hddd, 12'h999, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'h333, 12'h000, 12'h111, 12'h111, 12'h111, 12'h222, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h333, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hddd, 12'haaa, 12'h777, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h888, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h444, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hccc, 12'haaa, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h333, 12'h000, 12'h000, 12'h000, 12'h111, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hddd, 12'h999, 12'h555, 12'h777, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'h000, 12'h000, 12'h111, 12'h000, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hddd, 12'h999, 12'h666, 12'h999, 12'haaa, 12'hbbb, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h111, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hddd, 12'h999, 12'h999, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'haaa, 12'hccc, 12'h888, 12'h999, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h222, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h777, 12'h666, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h888, 12'h555, 12'h888, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h111, 12'h000, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h777, 12'h666, 12'haaa, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h000, 12'h000, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h333, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h777, 12'h777, 12'hccc, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'haaa, 12'h444, 12'h000, 12'h000, 12'h222, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h777, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h222, 12'h111, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h222, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h777, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h111, 12'h000, 12'h000, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 
12'h999, 12'haaa, 12'h777, 12'h777, 12'h999, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h555, 12'h111, 12'h000, 12'h333, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hbbb, 12'hccc, 12'h888, 12'h999, 12'hddd, 12'hbbb, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h222, 12'h000, 12'h111, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hddd, 12'hfff, 12'haaa, 12'h888, 12'hbbb, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h666, 12'h000, 12'h111, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 
12'hddd, 12'hfff, 12'haaa, 12'h999, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h111, 12'h000, 12'h111, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hddd, 12'heee, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h666, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h222, 12'h000, 12'h111, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h111, 12'h000, 12'h333, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h444, 12'h000, 12'h111, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h666, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h333, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h444, 12'h000, 12'h222, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h555, 12'h000, 12'h222, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'h777, 12'h444, 12'h444, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h555, 12'h444, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h444, 12'h111, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h333, 12'h000, 12'h333, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h444, 12'h000, 12'h222, 12'h999, 12'heee, 12'hddd, 12'heee, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'haaa, 12'h555, 12'h000, 12'h222, 12'h888, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'heee, 12'h777, 12'h666, 12'heee, 12'hfff, 12'hccc, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hccc, 12'hbbb, 12'hccc, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'h999, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h555, 12'h000, 12'h111, 12'h666, 12'hbbb, 12'hddd, 12'hccc, 12'hbbb, 12'heee, 12'h999, 12'h555, 12'hccc, 12'hddd, 12'hbbb, 12'hccc, 12'haaa, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h999, 12'hbbb, 12'h999, 12'h999, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'h777, 12'h777, 12'hbbb, 12'haaa, 12'haaa, 12'hbbb, 12'haaa, 12'h666, 12'h111, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'h999, 12'h777, 12'hccc, 12'h999, 12'h333, 12'h777, 12'h999, 12'haaa, 12'haaa, 12'h888, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h777, 12'h777, 12'h888, 12'h888, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'h999, 12'h444, 12'h111, 12'h333, 12'h444, 12'h555, 12'h666, 12'haaa, 12'hbbb, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h888, 12'h555, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h999, 12'h888, 12'h888, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'haaa, 12'h444, 12'h000, 12'h333, 12'h111, 12'h111, 12'h888, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'haaa, 12'h444, 12'h555, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hddd, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'haaa, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'haaa, 12'h222, 12'h222, 12'h666, 12'h666, 12'h666, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h555, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hddd, 12'hbbb, 12'h999, 12'h888, 12'h999, 12'h888, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h444, 12'h777, 12'h999, 12'h888, 12'h888, 12'h999, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'haaa, 12'h444, 12'h666, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 


// pipe 3, top to right 90 degrees

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h666, 12'h444, 12'haaa, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'h999, 12'h888, 12'h888, 12'h999, 12'h777, 12'h444, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h888, 12'h999, 12'h888, 12'h999, 12'hbbb, 12'hddd, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h666, 12'h666, 12'h666, 12'h222, 12'h222, 12'haaa, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hddd, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'h444, 12'haaa, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'h888, 12'h111, 12'h111, 12'h333, 12'h000, 12'h444, 12'haaa, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h999, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'h555, 12'h888, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hbbb, 12'haaa, 12'h666, 12'h555, 12'h444, 12'h333, 12'h111, 12'h444, 12'h999, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'hbbb, 12'haaa, 12'h888, 12'h888, 12'h777, 12'h777, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h999, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h888, 12'haaa, 12'haaa, 12'h999, 12'h777, 12'h333, 12'h999, 12'hccc, 12'h777, 12'h999, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h111, 12'h666, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'hbbb, 12'h777, 12'h777, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'h999, 12'h999, 12'hbbb, 12'h999, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'haaa, 12'hccc, 12'hbbb, 12'hddd, 12'hccc, 12'h555, 12'h999, 12'heee, 12'hbbb, 12'hccc, 12'hddd, 12'hbbb, 12'h666, 12'h111, 12'h000, 12'h555, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h999, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'hccc, 12'hbbb, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'hccc, 12'hfff, 12'heee, 12'h666, 12'h777, 12'heee, 12'hfff, 12'hddd, 12'hbbb, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h555, 12'haaa, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'heee, 12'hddd, 12'heee, 12'h999, 12'h222, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'h000, 12'h333, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h111, 12'h444, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h444, 12'h555, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h444, 12'h444, 12'h777, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h222, 12'h000, 12'h555, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h222, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'h000, 12'h222, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h666, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h111, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'h000, 12'h111, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h111, 12'h000, 12'h222, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h666, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'heee, 12'hddd, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h111, 12'h000, 12'h111, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'h999, 12'haaa, 12'hfff, 12'hddd, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h111, 12'h000, 12'h666, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 12'h888, 12'haaa, 12'hfff, 12'hddd, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h111, 12'h000, 12'h222, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'hbbb, 12'hddd, 12'h999, 12'h888, 12'hccc, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'h000, 12'h111, 12'h555, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h999, 12'h777, 12'h777, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h777, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h222, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h111, 12'h222, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h777, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'h000, 12'h000, 12'h444, 12'haaa, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hccc, 12'h777, 12'h777, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h333, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h000, 12'h000, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'haaa, 12'h666, 12'h777, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h000, 12'h111, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'h888, 12'h555, 12'h888, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h666, 12'h777, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h222, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'h999, 12'h888, 12'hccc, 12'haaa, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'h999, 12'h999, 12'hddd, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h000, 12'h111, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'hbbb, 12'haaa, 12'h999, 12'h666, 12'h999, 12'hddd, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'h000, 12'h111, 12'h000, 12'h000, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'h555, 12'h999, 12'hddd, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h111, 12'h000, 12'h000, 12'h000, 12'h333, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'haaa, 12'hccc, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'h888, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'haaa, 12'hddd, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h333, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h222, 12'h111, 12'h111, 12'h111, 12'h000, 12'h333, 12'h777, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'h999, 12'hddd, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h555, 12'h888, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'haaa, 12'hddd, 12'hbbb, 12'h999, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'h555, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'h444, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h333, 12'h555, 12'h777, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'haaa, 12'h777, 12'haaa, 12'hddd, 12'hccc, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h444, 12'h444, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'h999, 12'h555, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h444, 12'h444, 12'h444, 12'h555, 12'h666, 12'h666, 12'h555, 12'h888, 12'haaa, 12'h999, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h666, 12'h333, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h333, 12'h333, 12'h444, 12'h444, 12'h444, 12'h666, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h222, 12'h555, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h666, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h333, 12'h111, 12'h111, 12'h555, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h555, 12'h333, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h555, 12'h444, 12'h444, 12'h333, 12'h111, 12'h111, 12'h666, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'h444, 12'h444, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'haaa, 12'h777, 12'h111, 12'h000, 12'h000, 12'h666, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h444, 12'h555, 12'h777, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'hbbb, 12'hddd, 12'h999, 12'h000, 12'h000, 12'h111, 12'h555, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h666, 12'h444, 12'h444, 12'h666, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hccc, 12'h888, 12'h333, 12'h666, 12'h555, 12'h777, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h777, 12'h555, 12'h444, 12'h666, 12'h888, 12'haaa, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'h666, 12'hbbb, 12'heee, 12'hddd, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h666, 12'h444, 12'h444, 12'h555, 12'h777, 12'h888, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h666, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h888, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'haaa, 12'hccc, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h777, 12'h666, 12'h555, 12'h444, 12'h444, 12'h444, 12'h555, 12'h777, 12'hccc, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'h999, 12'h666, 12'hccc, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'hccc, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'hbbb, 12'hccc, 12'h999, 12'haaa, 12'heee, 12'hddd, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 12'h777, 12'h555, 12'h888, 12'h777, 12'h777, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h666, 12'h333, 12'h444, 12'h222, 12'h555, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h777, 12'h666, 12'h666, 12'h888, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hccc, 12'hddd, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 


// pipe four, bottom to right 90 degrees

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'h777, 12'h888, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h888, 12'h777, 12'h555, 12'h555, 12'h666, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h888, 12'h555, 12'h444, 12'h444, 12'h444, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'hccc, 12'haaa, 12'h888, 12'haaa, 12'hccc, 12'haaa, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'haaa, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'heee, 12'hccc, 12'h777, 12'h999, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h666, 12'h666, 12'h555, 12'h333, 12'h999, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h777, 12'h555, 12'h444, 12'h444, 12'h444, 12'h555, 12'h666, 12'h666, 12'h777, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h555, 12'h444, 12'h444, 12'h555, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hccc, 12'hbbb, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h888, 12'h555, 12'h444, 12'h444, 12'h666, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'haaa, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h666, 12'h444, 12'h444, 12'h777, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'h999, 12'h666, 12'h888, 12'haaa, 12'h999, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h666, 12'h444, 12'h555, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hddd, 12'hccc, 12'h555, 12'h111, 12'h666, 12'h888, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h555, 12'h222, 12'h555, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'haaa, 12'h444, 12'h111, 12'h666, 12'h888, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h333, 12'h444, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h666, 12'h555, 12'h333, 12'h333, 12'h666, 12'h999, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h444, 12'h333, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h777, 12'h555, 12'h333, 12'h222, 12'h222, 12'h111, 12'h000, 12'h111, 12'h000, 12'h222, 12'h777, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h222, 12'h555, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h777, 12'h444, 12'h333, 12'h222, 12'h222, 12'h444, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h444, 12'h222, 12'h444, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h333, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'h555, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'h555, 12'h444, 12'h333, 12'h444, 12'h555, 12'h555, 12'h666, 12'h999, 12'haaa, 12'haaa, 12'h888, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h444, 12'h444, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h777, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h444, 12'h555, 12'h777, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'haaa, 12'hbbb, 12'hddd, 12'heee, 12'hccc, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'h555, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h555, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h666, 12'h888, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hbbb, 12'hbbb, 12'hddd, 12'heee, 12'hccc, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h333, 12'h111, 12'h111, 12'h000, 12'h000, 12'h222, 12'h555, 12'h888, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h333, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h666, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h222, 12'h000, 12'h000, 12'h111, 12'h222, 12'h666, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h444, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h000, 12'h000, 12'h111, 12'h111, 12'h555, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h777, 12'haaa, 12'hddd, 12'hddd, 12'hbbb, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'h777, 12'h888, 12'hbbb, 12'hddd, 12'hbbb, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h000, 12'h111, 12'h000, 12'h444, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hddd, 12'hbbb, 12'h888, 12'hbbb, 12'hddd, 12'hbbb, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'haaa, 12'h777, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'haaa, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'h999, 12'h777, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h000, 12'h000, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'haaa, 12'hbbb, 12'haaa, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h333, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'h111, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hccc, 12'h999, 12'h888, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h111, 12'h111, 12'h000, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'heee, 12'haaa, 12'h777, 12'h999, 12'haaa, 12'h888, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h222, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h888, 12'haaa, 12'h999, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h000, 12'h000, 12'h000, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h777, 12'h888, 12'haaa, 12'h888, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h222, 12'h000, 12'h000, 12'h666, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'h999, 12'h777, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h111, 12'h000, 12'h333, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'hccc, 12'hbbb, 12'h888, 12'hbbb, 12'hddd, 12'hbbb, 12'haaa, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h222, 12'h111, 12'h111, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'hddd, 12'hfff, 12'hddd, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h000, 12'h111, 12'h444, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haaa, 12'hddd, 12'heee, 12'hccc, 12'hbbb, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h222, 12'h000, 12'h000, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'heee, 12'hddd, 12'hddd, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h000, 12'h000, 12'h333, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h222, 12'h000, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h111, 12'h000, 12'h222, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h333, 12'h000, 12'h000, 12'h555, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h111, 12'h000, 12'h222, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h000, 12'h000, 12'h333, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h111, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h000, 12'h333, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h000, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'heee, 12'hfff, 12'hbbb, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hccc, 12'h888, 12'h000, 12'h111, 12'h555, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'hccc, 12'heee, 12'hbbb, 12'h444, 12'haaa, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'h555, 12'h000, 12'h333, 12'h666, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'hbbb, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'hbbb, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hbbb, 12'hccc, 12'hbbb, 12'hbbb, 12'h999, 12'h555, 12'hccc, 12'hccc, 12'h888, 12'hccc, 12'hddd, 12'haaa, 12'h444, 12'h000, 12'h333, 12'h666, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'h777, 12'h999, 12'hddd, 12'hccc, 12'h999, 12'h888, 12'haaa, 12'hccc, 12'hddd, 12'hccc, 12'h999, 12'hddd, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'h777, 12'h999, 12'h888, 12'h777, 12'h666, 12'h777, 12'haaa, 12'h999, 12'h666, 12'h888, 12'h999, 12'h777, 12'h444, 12'h333, 12'h333, 12'h555, 12'h777, 12'h777, 12'h666, 12'h777, 12'h888, 12'h555, 12'h666, 12'h999, 12'h999, 12'h666, 12'h555, 12'h666, 12'h777, 12'h888, 12'h888, 12'h777, 12'h999, 12'h888, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h333, 12'h555, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h333, 12'h000, 12'h111, 12'h333, 12'h333, 12'h444, 12'h888, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h888, 12'h777, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'haaa, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'h444, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h000, 12'h000, 12'h111, 12'h111, 12'h444, 12'haaa, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h777, 12'hddd, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hddd, 12'h555, 12'h111, 12'h000, 12'h111, 12'h111, 12'h444, 12'h999, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h555, 12'h777, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h777, 12'h555, 12'h666, 12'h666, 12'h555, 12'h666, 12'h888, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 


//pipe five, left to top 90 degrees

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h888, 12'h666, 12'h555, 12'h666, 12'h666, 12'h555, 12'h777, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h777, 12'h555, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'h999, 12'h444, 12'h111, 12'h111, 12'h000, 12'h111, 12'h555, 12'hddd, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hddd, 12'h777, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'haaa, 12'h444, 12'h111, 12'h111, 12'h000, 12'h000, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'haaa, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h777, 12'h888, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h888, 12'h444, 12'h333, 12'h333, 12'h111, 12'h000, 12'h333, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h333, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h888, 12'h999, 12'h777, 12'h888, 12'h888, 12'h777, 12'h666, 12'h555, 12'h666, 12'h999, 12'h999, 12'h666, 12'h555, 12'h888, 12'h777, 12'h666, 12'h777, 12'h777, 12'h555, 12'h333, 12'h333, 12'h444, 12'h777, 12'h999, 12'h888, 12'h666, 12'h999, 12'haaa, 12'h777, 12'h666, 12'h777, 12'h888, 12'h999, 12'h777, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hddd, 12'h999, 12'hccc, 12'hddd, 12'hccc, 12'haaa, 12'h888, 12'h999, 12'hccc, 12'hddd, 12'h999, 12'h777, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h666, 12'h333, 12'h000, 12'h444, 12'haaa, 12'hddd, 12'hccc, 12'h888, 12'hccc, 12'hccc, 12'h555, 12'h999, 12'hbbb, 12'hbbb, 12'hccc, 12'hbbb, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'hbbb, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'hbbb, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h666, 12'h333, 12'h000, 12'h555, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'heee, 12'haaa, 12'h444, 12'hbbb, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h555, 12'h111, 12'h000, 12'h888, 12'hccc, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'hbbb, 12'hfff, 12'heee, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h444, 12'h000, 12'h000, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h444, 12'h000, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h444, 12'h000, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h333, 12'h000, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h111, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h111, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h555, 12'h000, 12'h000, 12'h333, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h222, 12'h000, 12'h111, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h222, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 
12'hddd, 12'heee, 12'hddd, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h000, 12'h000, 12'h222, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hccc, 12'heee, 12'hddd, 12'haaa, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h444, 12'h111, 12'h000, 12'h444, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hddd, 12'hfff, 12'hddd, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h111, 12'h111, 12'h222, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hbbb, 12'hddd, 12'hbbb, 12'h888, 12'hbbb, 12'hccc, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h333, 12'h000, 12'h111, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h999, 12'haaa, 12'h999, 12'h777, 12'h999, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h666, 12'h000, 12'h000, 12'h222, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h888, 12'haaa, 12'h888, 12'h777, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h000, 12'h000, 12'h000, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h999, 12'haaa, 12'h888, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h222, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h888, 12'haaa, 12'h999, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h111, 12'h111, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h999, 12'haaa, 12'haaa, 12'h888, 12'h999, 12'hccc, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h111, 12'h000, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'haaa, 12'hbbb, 12'haaa, 12'h888, 12'h999, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h000, 12'h000, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'haaa, 12'haaa, 12'h999, 12'h777, 12'h999, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'haaa, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h222, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'haaa, 12'hbbb, 12'haaa, 12'h777, 12'haaa, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h555, 12'h000, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hbbb, 12'hddd, 12'hbbb, 12'h888, 12'hbbb, 12'hddd, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h444, 12'h000, 12'h111, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hbbb, 12'hddd, 12'hbbb, 12'h888, 12'h777, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'hbbb, 12'hddd, 12'hddd, 12'haaa, 12'h777, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h555, 12'h111, 12'h111, 12'h000, 12'h000, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h444, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hccc, 12'hddd, 12'hddd, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h666, 12'h222, 12'h111, 12'h000, 12'h000, 12'h222, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h444, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 
12'hccc, 12'hddd, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h666, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h333, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 
12'hccc, 12'hddd, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h555, 12'h222, 12'h000, 12'h000, 12'h111, 12'h111, 12'h333, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 
12'hccc, 12'heee, 12'hddd, 12'hbbb, 12'hbbb, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h666, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h555, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h555, 12'h444, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'hccc, 12'heee, 12'hddd, 12'hbbb, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h777, 12'h555, 12'h444, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h777, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h444, 12'h444, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h888, 12'haaa, 12'haaa, 12'h999, 12'h666, 12'h555, 12'h555, 12'h444, 12'h333, 12'h444, 12'h555, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h555, 12'h888, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h333, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'h444, 12'h222, 12'h444, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h444, 12'h222, 12'h222, 12'h333, 12'h444, 12'h777, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h555, 12'h222, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 
12'h777, 12'h222, 12'h000, 12'h111, 12'h000, 12'h111, 12'h222, 12'h222, 12'h333, 12'h555, 12'h777, 12'h777, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h333, 12'h444, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 
12'h999, 12'h666, 12'h333, 12'h333, 12'h555, 12'h666, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h444, 12'h333, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'h888, 12'h666, 12'h111, 12'h444, 12'haaa, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h555, 12'h222, 12'h555, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'h888, 12'h666, 12'h111, 12'h555, 12'hccc, 12'hddd, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h555, 12'h444, 12'h666, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h999, 12'haaa, 12'h888, 12'h666, 12'h999, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h777, 12'h444, 12'h444, 12'h666, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'hfff, 12'haaa, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h666, 12'h444, 12'h444, 12'h555, 12'h888, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hccc, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'h555, 12'h444, 12'h444, 12'h555, 12'h777, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'h777, 12'h666, 12'h666, 12'h555, 12'h444, 12'h444, 12'h444, 12'h555, 12'h777, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'heee, 12'h999, 12'h333, 12'h555, 12'h666, 12'h666, 12'h777, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'heee, 12'h999, 12'h777, 12'hccc, 12'heee, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'heee, 12'haaa, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 
12'heee, 12'hfff, 12'heee, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'haaa, 12'hccc, 12'haaa, 12'h888, 12'haaa, 12'hccc, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h444, 12'h444, 12'h444, 12'h555, 12'h888, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 
12'h666, 12'h555, 12'h555, 12'h777, 12'h888, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 
12'h888, 12'h777, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 


// pipe 6, cross pipe

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h555, 12'h666, 12'h999, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hbbb, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h111, 12'h444, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h000, 12'h222, 12'h111, 12'h111, 12'h333, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'h666, 12'h666, 12'h666, 12'h333, 12'h333, 12'h333, 12'h777, 12'h999, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h999, 12'haaa, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'hccc, 12'hbbb, 12'hbbb, 12'h888, 12'h333, 12'h777, 12'haaa, 12'h999, 12'h666, 12'h999, 12'hbbb, 12'haaa, 12'h444, 12'h222, 12'h222, 12'h555, 12'h777, 12'h888, 12'h777, 12'h777, 12'h888, 12'h555, 12'h666, 12'haaa, 12'haaa, 12'h888, 12'h666, 12'h666, 12'h888, 12'haaa, 12'h999, 12'h777, 12'h999, 12'h999, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hddd, 12'hddd, 12'heee, 12'hccc, 12'h666, 12'h777, 12'hccc, 12'hccc, 12'haaa, 12'hccc, 12'heee, 12'hbbb, 12'h333, 12'h000, 12'h111, 12'h666, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'h888, 12'h999, 12'hccc, 12'hddd, 12'haaa, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'hddd, 12'haaa, 12'hbbb, 12'hccc, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hccc, 12'hfff, 12'hddd, 12'hbbb, 12'hccc, 12'hbbb, 12'h333, 12'h000, 12'h222, 12'h777, 12'hccc, 12'hddd, 12'hccc, 12'hddd, 12'hddd, 12'hbbb, 12'haaa, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'hfff, 12'heee, 12'h888, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hccc, 12'h444, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 
12'hbbb, 12'hbbb, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h111, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbbb, 12'hccc, 12'heee, 12'hbbb, 
12'h555, 12'h444, 12'h555, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h555, 12'h444, 12'h555, 12'hbbb, 12'haaa, 
12'h333, 12'h444, 12'h555, 12'h555, 12'h888, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h777, 12'h444, 12'h555, 12'h444, 12'h333, 12'haaa, 12'haaa, 
12'h666, 12'h888, 12'h888, 12'h666, 12'h999, 12'hbbb, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbbb, 12'h888, 12'h555, 12'h888, 12'h888, 12'h777, 12'hbbb, 12'hbbb, 
12'hbbb, 12'heee, 12'hddd, 12'h888, 12'haaa, 12'hccc, 12'h999, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'haaa, 12'hccc, 12'haaa, 12'h888, 12'heee, 12'heee, 12'hbbb, 12'hccc, 12'hbbb, 
12'hddd, 12'hfff, 12'hfff, 12'h999, 12'h999, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'h999, 12'haaa, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 
12'hccc, 12'hfff, 12'hfff, 12'h999, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h999, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 
12'hccc, 12'hfff, 12'hfff, 12'h888, 12'h444, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h777, 12'h333, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 
12'hccc, 12'hfff, 12'hfff, 12'h999, 12'h666, 12'h555, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h333, 12'h000, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'hddd, 12'h888, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h666, 12'h777, 12'haaa, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 
12'hccc, 12'hfff, 12'hfff, 12'haaa, 12'haaa, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'h777, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hddd, 12'haaa, 12'haaa, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 
12'hddd, 12'hfff, 12'hfff, 12'haaa, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'haaa, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hbbb, 
12'hbbb, 12'hddd, 12'hddd, 12'h888, 12'h666, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h666, 12'h999, 12'hddd, 12'hddd, 12'haaa, 12'hbbb, 12'haaa, 
12'h555, 12'h666, 12'h666, 12'h444, 12'haaa, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hccc, 12'h999, 12'h444, 12'h666, 12'h666, 12'h555, 12'hbbb, 12'haaa, 
12'h333, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hccc, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h888, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'hddd, 12'haaa, 12'h111, 12'h000, 12'h111, 12'h333, 12'hbbb, 12'haaa, 
12'h333, 12'h000, 12'h111, 12'h444, 12'h888, 12'haaa, 12'haaa, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h666, 12'h999, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h333, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'haaa, 
12'h333, 12'h000, 12'h111, 12'h444, 12'h333, 12'h444, 12'h555, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'haaa, 12'heee, 12'hddd, 12'h333, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h555, 12'h333, 12'h444, 12'h333, 12'h111, 12'h000, 12'h444, 12'hbbb, 12'haaa, 
12'h333, 12'h111, 12'h111, 12'h333, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'h999, 12'haaa, 12'h333, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h222, 12'h333, 12'h000, 12'h111, 12'h444, 12'hbbb, 12'haaa, 
12'h444, 12'h444, 12'h555, 12'h444, 12'h222, 12'h000, 12'h000, 12'h111, 12'h111, 12'h111, 12'h000, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h000, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h333, 12'h000, 12'h111, 12'h222, 12'h777, 12'hbbb, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h555, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h000, 12'h111, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h111, 12'h111, 12'h111, 12'h000, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h444, 12'h555, 12'h444, 12'h444, 12'hbbb, 12'hbbb, 
12'h888, 12'haaa, 12'haaa, 12'h666, 12'h555, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h777, 12'h777, 12'h555, 12'h777, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h777, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h555, 12'h777, 12'haaa, 12'haaa, 12'h888, 12'hbbb, 12'hbbb, 
12'haaa, 12'hddd, 12'hccc, 12'h888, 12'h777, 12'hbbb, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h777, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'h888, 12'hddd, 12'hddd, 12'haaa, 12'hbbb, 12'hbbb, 
12'haaa, 12'hccc, 12'hccc, 12'h777, 12'h888, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h777, 12'h888, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h777, 12'h888, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'haaa, 12'hccc, 12'hccc, 12'h777, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h444, 12'h333, 12'h666, 12'hbbb, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h888, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'haaa, 12'hccc, 12'hccc, 12'h777, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h333, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h888, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'haaa, 12'hccc, 12'hccc, 12'h777, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h111, 12'h111, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h888, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'haaa, 12'hccc, 12'hccc, 12'h777, 12'h555, 12'h888, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hddd, 12'heee, 12'hddd, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'h888, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'h888, 12'h555, 12'h888, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'haaa, 12'hccc, 12'hccc, 12'h777, 12'h777, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h777, 12'h777, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'haaa, 12'h777, 12'h888, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'haaa, 12'hccc, 12'hccc, 12'h777, 12'hbbb, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h111, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'h999, 12'h777, 12'h777, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hddd, 12'haaa, 12'h777, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'h999, 12'hbbb, 12'hbbb, 12'h666, 12'haaa, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h888, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'h888, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'h999, 12'h777, 12'hbbb, 12'hbbb, 12'h888, 12'hbbb, 12'hbbb, 
12'h777, 12'h999, 12'h999, 12'h666, 12'h777, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h666, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h666, 12'h666, 12'haaa, 12'h999, 12'h777, 12'hbbb, 12'hbbb, 
12'h888, 12'haaa, 12'h999, 12'h666, 12'h666, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'h777, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'h999, 12'h666, 12'h777, 12'haaa, 12'haaa, 12'h777, 12'hbbb, 12'hbbb, 
12'h888, 12'haaa, 12'h999, 12'h666, 12'h777, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'h666, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'hccc, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h777, 12'h666, 12'haaa, 12'haaa, 12'h777, 12'hbbb, 12'hbbb, 
12'h888, 12'haaa, 12'h999, 12'h666, 12'h999, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'haaa, 12'h333, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'hddd, 12'hbbb, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'h888, 12'h777, 12'haaa, 12'haaa, 12'h777, 12'hbbb, 12'haaa, 
12'h888, 12'haaa, 12'h999, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h777, 12'h999, 12'haaa, 12'h777, 12'hbbb, 12'haaa, 
12'h777, 12'h999, 12'h999, 12'h666, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h777, 12'h777, 12'h999, 12'h999, 12'h777, 12'hbbb, 12'hbbb, 
12'h888, 12'haaa, 12'h999, 12'h666, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h666, 12'haaa, 12'h999, 12'h777, 12'hbbb, 12'hbbb, 
12'haaa, 12'hddd, 12'hccc, 12'h777, 12'haaa, 12'hbbb, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'haaa, 12'hccc, 12'h999, 12'h777, 12'hccc, 12'hccc, 12'h999, 12'hbbb, 12'hbbb, 
12'hbbb, 12'hfff, 12'heee, 12'h777, 12'h999, 12'hbbb, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbbb, 12'h999, 12'h888, 12'heee, 12'heee, 12'hbbb, 12'hbbb, 12'hbbb, 
12'hbbb, 12'heee, 12'heee, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'heee, 12'heee, 12'hbbb, 12'hbbb, 12'hddd, 
12'hccc, 12'heee, 12'heee, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'heee, 12'heee, 12'hccc, 12'hddd, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h111, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'heee, 12'h999, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h333, 12'h000, 12'h111, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haaa, 12'heee, 12'heee, 12'h999, 12'h777, 12'hddd, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'h444, 12'h000, 12'h222, 12'h777, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'hccc, 12'hbbb, 12'hddd, 12'hddd, 12'h999, 12'h999, 12'hddd, 12'heee, 12'hccc, 12'hbbb, 12'hddd, 12'haaa, 12'h333, 12'h000, 12'h111, 12'h666, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'heee, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h888, 12'h999, 12'hbbb, 12'haaa, 12'h888, 12'hbbb, 12'hddd, 12'h999, 12'h333, 12'h222, 12'h111, 12'h555, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'h666, 12'h777, 12'hccc, 12'hccc, 12'h999, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'hbbb, 12'h999, 12'hbbb, 12'hccc, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h888, 12'h999, 12'haaa, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'h999, 12'h777, 12'h777, 12'h888, 12'h555, 12'h333, 12'h222, 12'h333, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h999, 12'h999, 12'h888, 12'h666, 12'h555, 12'h666, 12'h888, 12'h888, 12'h777, 12'h888, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h777, 12'h888, 12'hccc, 12'heee, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h222, 12'h222, 12'h333, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h888, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h666, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'h111, 12'h000, 12'h000, 12'h222, 12'haaa, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'heee, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'h666, 12'h999, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h666, 12'h111, 12'h222, 12'h222, 12'h222, 12'h333, 12'h999, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h888, 12'h999, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 

// pipe seven, blocked pipe

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h777, 12'h666, 12'h555, 12'h555, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h777, 12'h555, 12'h555, 12'h555, 12'h555, 12'h777, 12'h888, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h888, 12'h777, 12'h666, 12'h444, 12'h555, 12'h555, 12'h777, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h777, 12'h555, 12'h555, 12'h777, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'h999, 12'h777, 12'h555, 12'h444, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h666, 12'h444, 12'h666, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h666, 12'h555, 12'h666, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h555, 12'h444, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h444, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h444, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h444, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h888, 12'h555, 12'h333, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h555, 12'h888, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h666, 12'h555, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h444, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h444, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h555, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h555, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h000, 12'h111, 12'h222, 12'h333, 12'h000, 12'h000, 12'h111, 12'h222, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h555, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h111, 12'h000, 12'h000, 12'h333, 12'h444, 12'h444, 12'h666, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h666, 12'h444, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h000, 12'h111, 12'h000, 12'h000, 12'h444, 12'h777, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h666, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'h000, 12'h111, 12'h000, 12'h444, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h000, 12'h000, 12'h000, 12'h111, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'h000, 12'h000, 12'h000, 12'h111, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h111, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h444, 12'h111, 12'h111, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'h111, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'h000, 12'h000, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h111, 12'h000, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h111, 12'h000, 12'h000, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h111, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h444, 12'h000, 12'h111, 12'h555, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h555, 12'h000, 12'h000, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'h000, 12'h333, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h333, 12'h111, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h000, 12'h111, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h111, 12'h000, 12'h222, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h555, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h000, 12'h111, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h000, 12'h000, 12'h222, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h666, 12'h000, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h111, 12'h222, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h000, 12'h000, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'h111, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h555, 12'h000, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h222, 12'h333, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h000, 12'h000, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h111, 12'h222, 12'h333, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h333, 12'h333, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h111, 12'h666, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h666, 12'h222, 12'h111, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h111, 12'h000, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'h888, 12'h000, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'h000, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'h999, 12'h555, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h000, 12'h222, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hbbb, 12'h333, 12'h000, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h333, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'h333, 12'h000, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h111, 12'h000, 12'h555, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hccc, 12'haaa, 12'hfff, 12'hddd, 12'h444, 12'hccc, 12'hfff, 12'hddd, 12'hccc, 12'hbbb, 12'h000, 12'h111, 12'h666, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hbbb, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hddd, 12'hccc, 12'hddd, 12'hccc, 12'h555, 12'h000, 12'h111, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'hbbb, 12'h555, 12'hddd, 12'hfff, 12'haaa, 12'hddd, 12'hbbb, 
12'hbbb, 12'hddd, 12'heee, 12'hccc, 12'h555, 12'hddd, 12'hccc, 12'haaa, 12'hccc, 12'haaa, 12'h444, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'hccc, 12'hbbb, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hbbb, 12'hccc, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hccc, 12'hbbb, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'hddd, 12'hccc, 12'h999, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'h666, 12'h000, 12'h000, 12'h999, 12'hddd, 12'hbbb, 12'hddd, 12'hccc, 12'h555, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'hbbb, 
12'hbbb, 12'hccc, 12'hccc, 12'h999, 12'h777, 12'hbbb, 12'h777, 12'h999, 12'hbbb, 12'h777, 12'h777, 12'h333, 12'h555, 12'h888, 12'h777, 12'h888, 12'h777, 12'h666, 12'hbbb, 12'haaa, 12'h777, 12'h777, 12'h888, 12'hbbb, 12'h888, 12'haaa, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'haaa, 12'haaa, 12'h888, 12'hbbb, 12'h888, 12'h888, 12'h888, 12'haaa, 12'hccc, 12'h777, 12'h999, 12'h999, 12'h888, 12'h888, 12'h555, 12'h222, 12'h333, 12'h777, 12'hbbb, 12'h999, 12'h888, 12'hbbb, 12'h555, 12'h777, 12'haaa, 12'hbbb, 12'h999, 12'haaa, 
12'haaa, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'h777, 12'h333, 12'h555, 12'h888, 12'h444, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h888, 12'h999, 12'h999, 12'h888, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbbb, 12'h888, 12'h888, 12'h888, 12'h999, 12'h999, 12'h888, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'h888, 12'h444, 12'h444, 12'h333, 12'h333, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h777, 12'hccc, 
12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h888, 12'h999, 12'h777, 12'h666, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h555, 12'h555, 12'h555, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'haaa, 
12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h888, 12'h777, 12'h777, 12'h777, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h666, 12'h666, 12'h666, 12'h666, 12'h999, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'h999, 12'h666, 
12'h777, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'haaa, 12'h888, 12'h777, 12'h888, 12'h777, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'h888, 12'h888, 12'h888, 12'h999, 12'hbbb, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'haaa, 12'h888, 
12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h888, 12'h888, 12'h777, 12'h777, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'hddd, 12'h888, 12'h999, 12'haaa, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 
12'h666, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'h888, 12'h555, 12'h555, 12'h555, 12'h666, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hbbb, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'haaa, 12'hbbb, 12'hbbb, 12'haaa, 12'h666, 12'h999, 12'h777, 12'h666, 12'h999, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'haaa, 12'hbbb, 
12'h999, 12'hbbb, 12'haaa, 12'h777, 12'h555, 12'hbbb, 12'h888, 12'h999, 12'hccc, 12'h888, 12'h333, 12'h444, 12'h555, 12'h888, 12'h888, 12'haaa, 12'h999, 12'h888, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h888, 12'hbbb, 12'h888, 12'haaa, 12'haaa, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'hbbb, 12'h999, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'haaa, 12'hbbb, 12'h666, 12'h888, 12'h888, 12'h888, 12'h888, 12'h666, 12'h444, 12'h888, 12'h888, 12'hccc, 12'haaa, 12'h888, 12'hbbb, 12'h888, 12'haaa, 12'hccc, 12'hccc, 12'hbbb, 12'hddd, 
12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'h555, 12'hccc, 12'hddd, 12'hbbb, 12'hddd, 12'h999, 12'h111, 12'h111, 12'h666, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'h999, 12'hccc, 12'hddd, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hbbb, 12'hccc, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hbbb, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'hbbb, 12'hddd, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h222, 12'h444, 12'haaa, 12'hddd, 12'hbbb, 12'hccc, 12'hddd, 12'h555, 12'hccc, 12'heee, 12'hddd, 12'hbbb, 12'hfff, 
12'hddd, 12'haaa, 12'hfff, 12'hddd, 12'h555, 12'hbbb, 12'hfff, 12'hddd, 12'hbbb, 12'hccc, 12'h000, 12'h111, 12'h555, 12'hccc, 12'hddd, 12'hccc, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'hbbb, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h666, 12'h000, 12'h000, 12'hccc, 12'hccc, 12'hddd, 12'hfff, 12'hccc, 12'h444, 12'hddd, 12'hfff, 12'haaa, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h111, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h555, 12'h000, 12'h111, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h333, 12'h111, 12'h333, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h333, 12'h111, 12'h222, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'h333, 12'hbbb, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h111, 12'h111, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h555, 12'h999, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h000, 12'h000, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h111, 12'h000, 12'h888, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h111, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h111, 12'h222, 12'h666, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h666, 12'h000, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h444, 12'h333, 12'h333, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h333, 12'h222, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'h000, 12'h888, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h333, 12'h222, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h000, 12'h555, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h222, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h333, 12'h111, 12'h000, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h222, 12'h111, 12'h222, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h000, 12'h666, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hccc, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h000, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h111, 12'h000, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'h000, 12'h555, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h000, 12'h999, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h999, 12'h111, 12'h111, 12'h111, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h111, 12'h333, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h444, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h555, 12'h000, 12'h000, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h111, 12'h111, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h000, 12'h111, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h111, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h000, 12'h111, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h000, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h000, 12'h000, 12'h000, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'h000, 12'h000, 12'h777, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h777, 12'h000, 12'h111, 12'h000, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h111, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'haaa, 12'h444, 12'h000, 12'h111, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h000, 12'h000, 12'h000, 12'h777, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'h888, 12'h111, 12'h000, 12'h000, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h999, 12'h444, 12'h000, 12'h111, 12'h000, 12'h222, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h111, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'haaa, 12'h777, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h444, 12'h666, 12'h888, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h666, 12'h444, 12'h444, 12'h333, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h555, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h777, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h222, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h222, 12'h000, 12'h000, 12'h000, 12'h333, 12'h222, 12'h111, 12'h000, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h555, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h555, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h000, 12'h111, 12'h222, 12'h444, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h444, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h555, 12'h666, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h555, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h111, 12'h333, 12'h555, 12'h888, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'h444, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h777, 12'h444, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'h444, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h444, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h444, 12'h555, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h666, 12'h555, 12'h666, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h666, 12'h444, 12'h666, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h444, 12'h555, 12'h777, 12'h999, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h777, 12'h555, 12'h555, 12'h777, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h777, 12'h555, 12'h555, 12'h444, 12'h555, 12'h777, 12'h888, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'h999, 12'h999, 12'h888, 12'h777, 12'h666, 12'h555, 12'h555, 12'h555, 12'h777, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h777, 12'h666, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h555, 12'h555, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 


// starting point

12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'hbbb, 12'heee, 12'h999, 12'h000, 12'h444, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h222, 12'h444, 12'h000, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'h000, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h111, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h555, 12'h000, 12'h444, 12'h999, 12'h111, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h000, 12'h000, 12'h444, 12'haaa, 12'heee, 12'hfff, 12'h888, 12'h111, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h000, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h000, 12'h000, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h222, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'h222, 12'h999, 12'h999, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hbbb, 12'h000, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haaa, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h000, 12'h111, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h000, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h111, 12'h333, 12'hccc, 12'h999, 12'h111, 12'h000, 12'h222, 12'hbbb, 12'haaa, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h111, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h000, 12'haaa, 12'haaa, 12'h444, 12'h000, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'haaa, 12'h000, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h111, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h333, 12'h111, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h666, 12'heee, 12'haaa, 12'h000, 12'h000, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h111, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'haaa, 12'h777, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'h888, 12'h222, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h222, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'hddd, 12'heee, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'hddd, 12'hfff, 12'h888, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'h444, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h111, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'hddd, 12'hfff, 12'hddd, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h111, 12'h666, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h444, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'h555, 12'h222, 12'heee, 12'hfff, 12'haaa, 12'h000, 12'h222, 12'h111, 12'heee, 12'hbbb, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'haaa, 12'hfff, 12'h444, 12'h666, 12'h888, 12'h000, 12'h888, 12'h222, 12'h222, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h555, 12'h999, 12'h000, 12'hccc, 12'hddd, 12'h000, 12'h333, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h666, 12'h888, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'h111, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h111, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h000, 12'h777, 12'hfff, 12'hfff, 12'h555, 12'h222, 12'hccc, 12'hddd, 12'hbbb, 12'haaa, 12'h888, 12'h666, 12'h333, 12'h000, 12'h000, 12'h000, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h333, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'heee, 12'hfff, 12'haaa, 12'h000, 12'h888, 12'hfff, 12'heee, 12'heee, 12'h999, 12'h000, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h333, 12'h000, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h333, 12'h111, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'h000, 12'h222, 12'h111, 12'h111, 12'h222, 12'h222, 12'h111, 12'h000, 12'h000, 12'h222, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h111, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h333, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h999, 12'h777, 12'h000, 12'h555, 12'h999, 12'h999, 12'haaa, 12'hddd, 12'haaa, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'h444, 12'h333, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'h999, 12'h111, 12'hbbb, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'heee, 12'h333, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'h888, 12'h000, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'h999, 12'h777, 12'h000, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h333, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hddd, 12'h111, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h111, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h222, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h333, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h444, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h111, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h111, 12'h111, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h222, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h333, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h333, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h333, 12'h111, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h333, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h333, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h111, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h222, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h111, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h000, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h222, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 


// ending point


12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'haaa, 12'h888, 12'h555, 12'h333, 12'h111, 12'h111, 12'h000, 12'h111, 12'h000, 12'h111, 12'h666, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h444, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h333, 12'h222, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h666, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h222, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h666, 12'h666, 12'h888, 12'haaa, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'h222, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h666, 12'h666, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h333, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h666, 12'h555, 12'h777, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h555, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h555, 12'h666, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h888, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'h444, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h777, 12'h555, 12'h777, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'h777, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h666, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h888, 12'hccc, 12'h555, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h888, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'h777, 12'h444, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h666, 12'heee, 12'hccc, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h666, 12'hddd, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h444, 12'hddd, 12'hfff, 12'h888, 12'h111, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h222, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h333, 12'hddd, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'hccc, 12'hfff, 12'heee, 12'h444, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'hccc, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hccc, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h222, 12'hbbb, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h777, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hddd, 12'h666, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h222, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h111, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'h777, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h333, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'h999, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h888, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h666, 12'h111, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h222, 12'hccc, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'h999, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h111, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h444, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h555, 12'hddd, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h111, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h999, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h111, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h000, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h444, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h333, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h000, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h333, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h333, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h333, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'h999, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h888, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h777, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h111, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h111, 12'h999, 12'hfff, 12'heee, 12'h999, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h444, 12'h000, 12'h555, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h666, 12'haaa, 12'h888, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'hddd, 12'hfff, 12'heee, 12'haaa, 12'h444, 12'h111, 12'h555, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h333, 12'h666, 12'h777, 12'h444, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h777, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'haaa, 12'h888, 12'h555, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h222, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h555, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h333, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h111, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h777, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h111, 12'h999, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h444, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h777, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h666, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h888, 12'h666, 12'h777, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h888, 12'h777, 12'h777, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h999, 12'h888, 12'h999, 12'h999, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
};
	
reg [11:0] winning_screen [0:307200] = {12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haba, 12'haaa, 12'hbba, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hdee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hdde, 12'hccc, 12'hbbb, 12'habb, 12'hbbc, 12'hbbc, 12'hbcc, 12'hbcc, 12'hcdd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'h888, 12'h887, 12'h887, 12'h898, 12'h998, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h898, 12'h899, 12'h999, 12'h999, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hcdd, 12'hdee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hccd, 12'hbcc, 12'hbcc, 12'h9aa, 12'h889, 12'h788, 12'h788, 12'h778, 12'h778, 12'h788, 12'h788, 12'h899, 12'h99a, 12'habb, 12'hccc, 12'hcdd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h898, 12'h888, 12'h888, 12'h887, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h777, 12'h776, 12'h776, 12'h666, 12'h676, 12'h777, 12'h777, 12'h676, 12'h777, 12'h677, 12'h777, 12'h676, 12'h666, 12'h676, 12'h676, 12'h777, 12'h677, 12'h676, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hdde, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hcdd, 12'hbcc, 12'hbcc, 12'haab, 12'h899, 12'h899, 12'h788, 12'h667, 12'h567, 12'h677, 12'h667, 12'h566, 12'h566, 12'h566, 12'h567, 12'h566, 12'h566, 12'h788, 12'h899, 12'h9aa, 12'haab, 12'hbbc, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h999, 12'h888, 12'h888, 12'h787, 12'h787, 12'h777, 12'h676, 12'h776, 12'h776, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h655, 12'h665, 12'h565, 12'h565, 12'h565, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'habb, 12'hcdd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbcc, 12'haab, 12'h9aa, 12'h899, 12'h778, 12'h667, 12'h567, 12'h566, 12'h456, 12'h456, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h566, 12'h677, 12'h678, 12'h788, 12'h889, 12'h999, 12'habb, 12'hccc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heff, 12'heff, 12'heff, 12'heff, 12'heef, 12'heff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbba, 12'haaa, 12'h999, 12'h999, 12'h898, 12'h888, 12'h888, 12'h787, 12'h777, 12'h777, 12'h666, 12'h665, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h565, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h665, 12'h565, 12'h565, 12'h666, 12'h666, 12'h566, 12'h566, 12'h666, 12'h566, 12'h666, 12'h666, 12'h677, 12'h777, 12'h899, 12'habb, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'haaa, 12'h9aa, 12'h899, 12'h788, 12'h677, 12'h566, 12'h566, 12'h566, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h678, 12'h788, 12'h889, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 
12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h666, 12'h665, 12'h665, 12'h565, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h565, 12'h555, 12'h555, 12'h665, 12'h666, 12'h665, 12'h565, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h777, 12'h9aa, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'h889, 12'h788, 12'h677, 12'h567, 12'h566, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h355, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h566, 12'h788, 12'h9aa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heff, 12'heee, 12'hdee, 12'hdee, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'heee, 12'hdee, 12'hdde, 12'hddd, 
12'hdee, 12'heee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'haaa, 12'haaa, 12'haa9, 12'h999, 12'h998, 12'h888, 12'h887, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h666, 12'h666, 12'h565, 12'h555, 12'h555, 12'h665, 12'h665, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h777, 12'h999, 12'hbcc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h999, 12'h677, 12'h677, 12'h566, 12'h556, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h355, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h889, 12'haaa, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hcdd, 12'hccc, 12'hccd, 12'hcdd, 12'hddd, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hcdd, 12'hccd, 12'hccc, 
12'hcdd, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heed, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h999, 12'h999, 12'h888, 12'h888, 12'h887, 12'h777, 12'h777, 12'h776, 12'h676, 12'h676, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h666, 12'h665, 12'h665, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h565, 12'h565, 12'h555, 12'h555, 12'h555, 12'h665, 12'h665, 12'h665, 12'h666, 12'h665, 12'h665, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h555, 12'h555, 12'h566, 12'h666, 12'h777, 12'h777, 12'h788, 12'h9aa, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h999, 12'h788, 12'h778, 12'h777, 12'h677, 12'h677, 12'h677, 12'h566, 12'h566, 12'h556, 12'h455, 12'h455, 12'h345, 12'h345, 12'h455, 12'h355, 12'h355, 12'h355, 12'h345, 12'h455, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h566, 12'h677, 12'h889, 12'hccd, 12'heee, 12'heef, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdee, 12'hdee, 12'hddd, 12'hcdd, 12'hbcc, 12'habb, 12'hbbb, 12'hccc, 12'hccd, 12'hccd, 12'hccd, 12'hccc, 12'hccc, 12'hccd, 12'hccd, 12'hbcc, 12'hbbc, 12'hbbb, 
12'hbcc, 12'hccc, 12'hcdd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heff, 12'heff, 12'heff, 12'heff, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hddd, 12'hbbb, 12'hbba, 12'haaa, 12'haaa, 12'h999, 12'h998, 12'h888, 12'h888, 12'h777, 12'h777, 12'h776, 12'h776, 12'h777, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h555, 12'h665, 12'h665, 12'h665, 12'h655, 12'h655, 12'h555, 12'h555, 12'h555, 12'h565, 12'h555, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h777, 12'h788, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haab, 12'h788, 12'h677, 12'h566, 12'h566, 12'h566, 12'h456, 12'h455, 12'h456, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h355, 12'h345, 12'h344, 12'h344, 12'h345, 12'h345, 12'h455, 12'h455, 12'h355, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h455, 12'h456, 12'h456, 12'h566, 12'h999, 12'hbcc, 12'hdee, 12'heee, 12'heff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hddd, 12'hddd, 12'hcdd, 12'hcdd, 12'hccd, 12'hbbc, 12'h9aa, 12'h9aa, 12'hbbb, 12'hbbb, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hbcc, 12'habb, 12'haab, 12'h9aa, 
12'habb, 12'hbbc, 12'hbcc, 12'hccd, 12'hccc, 12'hccd, 12'hcdd, 12'hcdd, 12'hccd, 12'hccd, 12'hddd, 12'hdde, 12'hdee, 12'heef, 12'heef, 12'heef, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 
12'hbbb, 12'hbba, 12'haaa, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h887, 12'h777, 12'h777, 12'h776, 12'h676, 12'h776, 12'h776, 12'h666, 12'h665, 12'h665, 12'h665, 12'h655, 12'h655, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h555, 12'h555, 12'h665, 12'h665, 12'h555, 12'h555, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h565, 12'h565, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h565, 12'h666, 12'h555, 12'h555, 12'h666, 12'h677, 12'h788, 12'h777, 12'h788, 12'h9aa, 12'hbbb, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hbcc, 12'h999, 12'h677, 12'h677, 12'h566, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h355, 12'h345, 12'h345, 12'h344, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h456, 12'h456, 12'h556, 12'h567, 12'h99a, 12'hccc, 12'hdde, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hddd, 12'hbcc, 12'hbcc, 12'hccd, 12'hccd, 12'hccd, 12'hbbb, 12'h99a, 12'h899, 12'haaa, 12'haaa, 12'h9aa, 12'haaa, 12'habb, 12'habb, 12'hbbb, 12'habb, 12'h9aa, 12'h99a, 12'h899, 
12'h9aa, 12'haab, 12'habb, 12'habb, 12'habb, 12'hbcc, 12'hccd, 12'hbbc, 12'haab, 12'hbbc, 12'hbcc, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hddd, 12'hbbb, 
12'hbba, 12'haaa, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h887, 12'h777, 12'h776, 12'h776, 12'h776, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h655, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h655, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h555, 12'h565, 12'h666, 12'h666, 12'h666, 12'h899, 12'haaa, 12'hbcc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h899, 12'h777, 12'h566, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h355, 12'h355, 12'h345, 12'h344, 12'h345, 12'h355, 12'h455, 12'h455, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h677, 12'h999, 
12'hccc, 12'hdee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'haab, 12'haab, 12'hccc, 12'hbcc, 12'hbbc, 12'haab, 12'h9aa, 12'h788, 12'h9aa, 12'h9aa, 12'h888, 12'h888, 12'h9aa, 12'haab, 12'haab, 12'h9aa, 12'h9aa, 12'h99a, 12'h889, 
12'h99a, 12'h9aa, 12'h9aa, 12'h9aa, 12'h9ab, 12'habb, 12'habb, 12'h99a, 12'h899, 12'habb, 12'habc, 12'hbbc, 12'hccd, 12'hccd, 12'hcdd, 12'hccd, 12'hccd, 12'hccd, 12'hcdd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 
12'haaa, 12'haa9, 12'h999, 12'h888, 12'h888, 12'h887, 12'h777, 12'h777, 12'h666, 12'h676, 12'h776, 12'h776, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h655, 12'h666, 12'h666, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h665, 12'h565, 12'h665, 12'h665, 12'h565, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h565, 12'h565, 12'h565, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h888, 12'h999, 12'hccc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hcdd, 12'hbcc, 12'h99a, 12'h677, 12'h677, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h345, 12'h445, 12'h345, 12'h445, 12'h345, 12'h345, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h566, 12'h567, 12'h677, 
12'h899, 12'hbbb, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccc, 12'hbbb, 12'haaa, 12'h9aa, 12'hbbb, 12'hbbc, 12'hbbb, 12'haaa, 12'h9aa, 12'h788, 12'h899, 12'h99a, 12'h778, 12'h677, 12'h788, 12'h999, 12'h99a, 12'h999, 12'haaa, 12'h99a, 12'h788, 
12'h899, 12'h899, 12'h889, 12'h99a, 12'h9aa, 12'haab, 12'h99a, 12'h788, 12'h89a, 12'haab, 12'habb, 12'hbcc, 12'hbcc, 12'hbbc, 12'habc, 12'habb, 12'habc, 12'habc, 12'hbcc, 12'hcdd, 12'hdde, 12'hdee, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 
12'haa9, 12'h999, 12'h998, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h766, 12'h776, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h655, 12'h565, 12'h565, 12'h565, 12'h555, 12'h565, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h777, 12'h999, 12'hccc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbcc, 12'haaa, 12'h777, 12'h778, 12'h667, 12'h456, 12'h556, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h355, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h455, 12'h345, 12'h345, 12'h455, 12'h445, 12'h445, 12'h345, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h566, 12'h566, 12'h567, 
12'h778, 12'h899, 12'habb, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hccc, 12'haaa, 12'h9aa, 12'h99a, 12'h9aa, 12'habb, 12'hbbc, 12'h9aa, 12'h9aa, 12'h888, 12'h788, 12'h999, 12'h788, 12'h777, 12'h778, 12'h778, 12'h778, 12'h888, 12'h899, 12'h899, 12'h888, 
12'h888, 12'h778, 12'h778, 12'h889, 12'h99a, 12'haab, 12'h788, 12'h778, 12'h9aa, 12'haab, 12'habb, 12'hbbc, 12'haab, 12'h89a, 12'h789, 12'h9aa, 12'haab, 12'h9ab, 12'hbbc, 12'hccd, 12'hcdd, 12'hcdd, 12'hccd, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbba, 12'haaa, 12'haa9, 
12'h999, 12'h998, 12'h888, 12'h887, 12'h777, 12'h777, 12'h776, 12'h666, 12'h666, 12'h776, 12'h776, 12'h666, 12'h666, 12'h776, 12'h666, 12'h665, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h665, 12'h565, 12'h555, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h454, 12'h554, 12'h555, 12'h555, 12'h666, 12'h676, 12'h677, 12'h777, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h889, 12'h788, 12'h677, 12'h566, 12'h456, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h445, 12'h345, 12'h445, 12'h445, 12'h456, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h355, 12'h456, 12'h456, 12'h566, 
12'h567, 12'h677, 12'h889, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'haaa, 12'h999, 12'h999, 12'h888, 12'h99a, 12'hbbb, 12'haaa, 12'h99a, 12'h889, 12'h788, 12'h889, 12'h889, 12'h777, 12'h788, 12'h777, 12'h667, 12'h667, 12'h777, 12'h778, 12'h778, 
12'h778, 12'h777, 12'h777, 12'h788, 12'h99a, 12'h99a, 12'h677, 12'h899, 12'haab, 12'haaa, 12'h9aa, 12'habb, 12'h899, 12'h778, 12'h789, 12'h9aa, 12'h9aa, 12'h9aa, 12'haab, 12'habb, 12'h9ab, 12'h899, 12'h99a, 12'habb, 12'hbbc, 12'hbbc, 12'hbbc, 12'habb, 12'habb, 12'hbbc, 12'hccd, 12'hcdd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haaa, 12'haaa, 12'haa9, 12'h999, 
12'h999, 12'h888, 12'h888, 12'h888, 12'h776, 12'h666, 12'h666, 12'h666, 12'h766, 12'h776, 12'h777, 12'h776, 12'h777, 12'h777, 12'h666, 12'h666, 12'h665, 12'h665, 12'h555, 12'h555, 12'h655, 12'h555, 12'h555, 12'h665, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h565, 12'h666, 12'h666, 12'h666, 12'h888, 12'haaa, 12'hcdd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h9aa, 12'h455, 12'h355, 12'h556, 12'h566, 12'h566, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h345, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h344, 12'h345, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h445, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 
12'h456, 12'h556, 12'h567, 12'h778, 12'h99a, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hcdd, 12'habb, 12'h888, 12'h788, 12'h778, 12'h888, 12'haaa, 12'haab, 12'h99a, 12'h899, 12'h889, 12'h889, 12'h888, 12'h778, 12'h778, 12'h777, 12'h667, 12'h666, 12'h667, 12'h667, 12'h677, 
12'h677, 12'h677, 12'h677, 12'h888, 12'h999, 12'h888, 12'h778, 12'h999, 12'h99a, 12'haaa, 12'haab, 12'h999, 12'h788, 12'h778, 12'h889, 12'h889, 12'h99a, 12'h899, 12'h789, 12'h788, 12'h788, 12'h789, 12'h99a, 12'h9aa, 12'h899, 12'h788, 12'h778, 12'h788, 12'h899, 12'haab, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haaa, 12'haa9, 12'h998, 12'h998, 12'h998, 
12'h888, 12'h887, 12'h887, 12'h887, 12'h776, 12'h665, 12'h665, 12'h666, 12'h666, 12'h766, 12'h776, 12'h777, 12'h777, 12'h777, 12'h766, 12'h665, 12'h665, 12'h555, 12'h555, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h565, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h655, 12'h665, 12'h555, 12'h554, 12'h665, 12'h665, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h554, 12'h544, 12'h554, 12'h554, 12'h454, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h777, 12'h999, 12'hbbb, 12'hdde, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbcc, 12'h566, 12'h355, 12'h345, 12'h345, 12'h345, 12'h566, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h345, 12'h455, 12'h445, 12'h344, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h344, 12'h344, 12'h345, 12'h344, 12'h344, 12'h344, 12'h455, 12'h445, 12'h455, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h445, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 
12'h456, 12'h456, 12'h566, 12'h566, 12'h778, 12'hbbc, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hccc, 12'hbbc, 12'h889, 12'h677, 12'h777, 12'h777, 12'h889, 12'haaa, 12'h9aa, 12'h888, 12'h888, 12'h899, 12'h788, 12'h777, 12'h777, 12'h777, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h777, 12'h777, 12'h888, 12'h889, 12'h99a, 12'h889, 12'h788, 12'h777, 12'h788, 12'h777, 12'h778, 12'h889, 12'h788, 12'h678, 12'h678, 12'h899, 12'h99a, 12'h788, 12'h778, 12'h677, 12'h667, 12'h678, 12'h778, 12'h889, 12'h99a, 12'h889, 12'h899, 12'h9aa, 12'haab, 12'hbcc, 12'hddd, 12'hdee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdc, 12'hbbb, 12'haaa, 12'haa9, 12'h999, 12'h888, 12'h888, 12'h888, 
12'h887, 12'h777, 12'h776, 12'h777, 12'h666, 12'h665, 12'h655, 12'h665, 12'h666, 12'h666, 12'h776, 12'h776, 12'h776, 12'h777, 12'h776, 12'h666, 12'h655, 12'h555, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h665, 12'h554, 12'h554, 12'h554, 12'h665, 12'h665, 12'h555, 12'h665, 12'h666, 12'h665, 12'h554, 12'h554, 12'h544, 12'h444, 12'h544, 12'h555, 12'h555, 12'h554, 12'h544, 12'h554, 12'h554, 12'h454, 12'h554, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h777, 12'h888, 12'habb, 12'hdee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbc, 12'h888, 12'h455, 12'h355, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h345, 12'h445, 12'h445, 12'h345, 12'h344, 12'h344, 12'h445, 12'h345, 12'h344, 12'h334, 12'h345, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 12'h445, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 
12'h455, 12'h455, 12'h455, 12'h556, 12'h567, 12'h889, 12'hbbb, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hccc, 12'hbcc, 12'h999, 12'h788, 12'h677, 12'h677, 12'h778, 12'h999, 12'h9aa, 12'h888, 12'h788, 12'h899, 12'h888, 12'h666, 12'h777, 12'h777, 12'h777, 12'h667, 12'h666, 12'h667, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h888, 12'h788, 12'h777, 12'h666, 12'h777, 12'h888, 12'h777, 12'h777, 12'h778, 12'h677, 12'h777, 12'h788, 12'h889, 12'h788, 12'h677, 12'h667, 12'h677, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h889, 12'h9aa, 12'hbbc, 12'hccd, 12'hdde, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbba, 12'haaa, 12'haa9, 12'h999, 12'h888, 12'h877, 12'h887, 12'h887, 
12'h887, 12'h777, 12'h776, 12'h766, 12'h666, 12'h665, 12'h555, 12'h665, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h777, 12'h776, 12'h766, 12'h655, 12'h555, 12'h665, 12'h666, 12'h666, 12'h665, 12'h565, 12'h554, 12'h655, 12'h555, 12'h665, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h666, 12'h666, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h544, 12'h554, 12'h554, 12'h444, 12'h444, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h776, 12'h777, 12'haaa, 12'hcdd, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h677, 12'h566, 12'h455, 12'h355, 12'h355, 12'h345, 12'h345, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h344, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h445, 12'h345, 12'h345, 12'h344, 12'h445, 12'h445, 12'h344, 12'h344, 12'h445, 12'h345, 12'h345, 12'h445, 12'h345, 12'h445, 12'h445, 12'h445, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 
12'h455, 12'h455, 12'h455, 12'h455, 12'h566, 12'h667, 12'h778, 12'habb, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbbb, 12'hbbb, 12'h9aa, 12'h888, 12'h778, 12'h677, 12'h677, 12'h788, 12'h999, 12'h999, 12'h788, 12'h888, 12'h999, 12'h777, 12'h666, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h788, 12'h888, 12'h677, 12'h777, 12'h667, 12'h666, 12'h777, 12'h778, 12'h677, 12'h667, 12'h667, 12'h667, 12'h777, 12'h777, 12'h777, 12'h667, 12'h667, 12'h677, 12'h778, 12'h889, 12'h889, 12'h9aa, 12'hbbc, 12'hbbc, 12'hbcc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 
12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbba, 12'haaa, 12'haaa, 12'h999, 12'h888, 12'h887, 12'h776, 12'h887, 12'h887, 
12'h777, 12'h777, 12'h776, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h655, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h655, 12'h555, 12'h666, 12'h766, 12'h776, 12'h665, 12'h555, 12'h554, 12'h555, 12'h554, 12'h554, 12'h544, 12'h554, 12'h554, 12'h554, 12'h555, 12'h665, 12'h665, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h554, 12'h554, 12'h544, 12'h554, 12'h554, 12'h554, 12'h444, 12'h454, 12'h554, 12'h554, 12'h454, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h999, 12'hccc, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h778, 12'h566, 12'h455, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h345, 12'h344, 12'h344, 12'h344, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h345, 12'h455, 12'h345, 12'h345, 12'h455, 12'h345, 12'h344, 12'h345, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 
12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h556, 12'h566, 12'h788, 12'hcdd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'habb, 12'h9aa, 12'h999, 12'h889, 12'h778, 12'h777, 12'h667, 12'h777, 12'h888, 12'h889, 12'h888, 12'h778, 12'h889, 12'h888, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h676, 12'h676, 12'h777, 12'h777, 12'h666, 12'h888, 12'h777, 12'h666, 12'h667, 12'h666, 12'h677, 12'h777, 12'h777, 12'h666, 12'h666, 12'h667, 12'h667, 12'h767, 12'h767, 12'h667, 12'h667, 12'h667, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h788, 12'h788, 12'h889, 12'h99a, 12'habb, 12'hccc, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccb, 12'hbba, 12'haaa, 12'haa9, 12'h999, 12'h888, 12'h777, 12'h777, 12'h777, 12'h888, 12'h887, 
12'h777, 12'h777, 12'h776, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h555, 12'h655, 12'h666, 12'h665, 12'h666, 12'h666, 12'h665, 12'h665, 12'h555, 12'h655, 12'h666, 12'h776, 12'h666, 12'h555, 12'h554, 12'h555, 12'h554, 12'h554, 12'h444, 12'h444, 12'h554, 12'h554, 12'h554, 12'h555, 12'h665, 12'h655, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h443, 12'h544, 12'h444, 12'h454, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h454, 12'h565, 12'h666, 12'h666, 12'h777, 12'h999, 12'hbcc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h9aa, 12'h566, 12'h455, 12'h355, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h445, 12'h445, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 
12'h455, 12'h455, 12'h455, 12'h556, 12'h456, 12'h456, 12'h456, 12'h567, 12'h99a, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haab, 12'h999, 12'h888, 12'h889, 12'h788, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h788, 12'h778, 12'h888, 12'h888, 12'h777, 12'h666, 12'h666, 12'h666, 12'h776, 12'h766, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h888, 12'h777, 12'h666, 12'h666, 12'h666, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h767, 12'h767, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h777, 12'h788, 12'h899, 12'haaa, 12'hbbb, 12'hbbc, 12'hccd, 12'hdee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haab, 12'habb, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hddd, 
12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h999, 12'h898, 12'h888, 12'h777, 12'h776, 12'h776, 12'h887, 12'h777, 
12'h776, 12'h776, 12'h666, 12'h666, 12'h655, 12'h665, 12'h666, 12'h666, 12'h555, 12'h665, 12'h665, 12'h655, 12'h665, 12'h655, 12'h665, 12'h665, 12'h555, 12'h665, 12'h665, 12'h666, 12'h665, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h443, 12'h544, 12'h554, 12'h555, 12'h555, 12'h555, 12'h665, 12'h554, 12'h544, 12'h554, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h443, 12'h444, 12'h554, 12'h544, 12'h544, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hcdd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h889, 12'h677, 12'h455, 12'h355, 12'h345, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h345, 12'h344, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h345, 12'h344, 12'h345, 12'h455, 12'h345, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h345, 12'h455, 12'h345, 12'h345, 
12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h566, 12'h99a, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdee, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h888, 12'h777, 12'h777, 12'h667, 12'h667, 12'h777, 12'h777, 12'h878, 12'h888, 12'h888, 12'h888, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h767, 12'h667, 12'h667, 12'h777, 12'h778, 12'h788, 12'h788, 12'h888, 12'h889, 12'h899, 12'h99a, 12'haab, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'haaa, 12'h9aa, 12'h999, 12'h999, 12'h999, 12'h899, 12'h899, 12'h999, 12'h999, 12'h999, 12'h99a, 12'h9aa, 12'haaa, 12'haaa, 12'haab, 12'habb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbc, 
12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haaa, 12'h999, 12'h998, 12'h888, 12'h887, 12'h777, 12'h766, 12'h666, 12'h766, 12'h877, 12'h777, 
12'h776, 12'h776, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h665, 12'h655, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h554, 12'h555, 12'h555, 12'h655, 12'h666, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h444, 12'h443, 12'h443, 12'h554, 12'h655, 12'h655, 12'h555, 12'h555, 12'h554, 12'h544, 12'h554, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h544, 12'h554, 12'h444, 12'h443, 12'h444, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h565, 12'h565, 12'h566, 12'h566, 12'h677, 12'h777, 12'h999, 12'hbcc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'h99a, 12'h788, 12'h566, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h355, 12'h455, 12'h455, 12'h455, 12'h344, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 
12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h566, 12'h677, 12'haaa, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767, 12'h767, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h777, 12'h778, 12'h888, 12'h899, 12'h9aa, 12'habb, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hbcc, 12'hbbb, 12'habb, 12'haaa, 12'haaa, 12'h99a, 12'h999, 12'h999, 12'h899, 12'h899, 12'h889, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h889, 12'h889, 12'h889, 12'h889, 12'h889, 12'h999, 12'h999, 12'h99a, 12'h9aa, 12'h9aa, 12'haaa, 12'haab, 
12'hbbb, 12'hbbc, 12'hccc, 12'hcdd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddc, 12'hbbb, 12'h999, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h666, 12'h665, 12'h776, 12'h777, 12'h776, 
12'h776, 12'h666, 12'h665, 12'h555, 12'h665, 12'h666, 12'h666, 12'h665, 12'h655, 12'h555, 12'h554, 12'h554, 12'h555, 12'h655, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h655, 12'h444, 12'h544, 12'h554, 12'h554, 12'h444, 12'h444, 12'h554, 12'h554, 12'h555, 12'h555, 12'h655, 12'h655, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h444, 12'h444, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h565, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h888, 12'h888, 12'hbbb, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbc, 12'h778, 12'h667, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h345, 12'h344, 12'h345, 12'h344, 12'h345, 
12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h566, 12'h788, 12'hbcc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767, 12'h766, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h777, 12'h777, 12'h778, 12'h888, 12'h999, 12'haaa, 12'hbbc, 12'hcdd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'h99a, 12'h99a, 12'h899, 12'h889, 12'h889, 12'h788, 12'h788, 12'h788, 12'h788, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h788, 12'h889, 12'h889, 12'h889, 12'h889, 12'h899, 12'h899, 12'h899, 12'h999, 12'h9aa, 
12'haaa, 12'haab, 12'hbbb, 12'hccc, 12'hccd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haa9, 12'h888, 12'h887, 12'h887, 12'h777, 12'h776, 12'h766, 12'h665, 12'h665, 12'h777, 12'h776, 12'h666, 
12'h666, 12'h665, 12'h555, 12'h555, 12'h666, 12'h777, 12'h666, 12'h665, 12'h555, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h544, 12'h554, 12'h555, 12'h555, 12'h544, 12'h444, 12'h544, 12'h554, 12'h444, 12'h444, 12'h554, 12'h554, 12'h544, 12'h544, 12'h555, 12'h655, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h544, 12'h444, 12'h554, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h565, 12'h666, 12'h666, 12'h666, 12'h566, 12'h777, 12'h888, 12'haaa, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h667, 12'h566, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h345, 12'h345, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h244, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h445, 12'h345, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 
12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h556, 12'h778, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h99a, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h777, 12'h778, 12'h889, 12'h99a, 12'hbbb, 12'hccd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hcdd, 12'hccc, 12'hccc, 12'hbbc, 12'hbbb, 12'haab, 12'haab, 12'h9aa, 12'h99a, 12'h99a, 12'h89a, 12'h889, 12'h789, 12'h788, 12'h778, 12'h778, 12'h788, 12'h778, 12'h778, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h678, 12'h788, 12'h788, 12'h788, 12'h788, 12'h889, 12'h889, 12'h889, 12'h889, 12'h899, 
12'h99a, 12'h99a, 12'haaa, 12'hbbb, 12'hbbc, 12'hccc, 12'hcdd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'haa9, 12'h998, 12'h888, 12'h777, 12'h777, 12'h776, 12'h666, 12'h666, 12'h665, 12'h665, 12'h776, 12'h666, 12'h666, 
12'h665, 12'h555, 12'h554, 12'h555, 12'h776, 12'h887, 12'h666, 12'h655, 12'h555, 12'h554, 12'h555, 12'h554, 12'h554, 12'h555, 12'h555, 12'h554, 12'h544, 12'h554, 12'h554, 12'h554, 12'h544, 12'h544, 12'h554, 12'h544, 12'h444, 12'h554, 12'h554, 12'h554, 12'h543, 12'h554, 12'h655, 12'h655, 12'h554, 12'h554, 12'h544, 12'h544, 12'h444, 12'h554, 12'h554, 12'h554, 12'h554, 12'h444, 12'h554, 12'h554, 12'h554, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'habb, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbcc, 12'h788, 12'h566, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h455, 12'h445, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h455, 12'h455, 12'h345, 12'h345, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h445, 12'h345, 12'h345, 12'h445, 12'h355, 12'h345, 12'h345, 12'h345, 
12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h889, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h888, 12'h878, 12'h777, 12'h777, 12'h766, 12'h767, 12'h766, 12'h777, 12'h777, 12'h766, 12'h767, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h777, 12'h778, 12'h888, 12'h99a, 12'habb, 12'hccd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'habb, 12'haab, 12'haab, 12'h9aa, 12'h99a, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h789, 12'h778, 12'h778, 12'h678, 12'h778, 12'h678, 12'h677, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h678, 12'h788, 12'h788, 12'h789, 12'h789, 12'h788, 12'h788, 12'h889, 12'h889, 
12'h889, 12'h899, 12'h99a, 12'haaa, 12'haab, 12'hbbb, 12'hbcc, 12'hccc, 12'hccd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h999, 12'h888, 12'h887, 12'h777, 12'h776, 12'h776, 12'h776, 12'h666, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h555, 12'h554, 12'h554, 12'h555, 12'h776, 12'h776, 12'h665, 12'h665, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h544, 12'h544, 12'h444, 12'h444, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h554, 12'h544, 12'h554, 12'h544, 12'h544, 12'h544, 12'h554, 12'h544, 12'h554, 12'h444, 12'h444, 12'h554, 12'h444, 12'h554, 12'h554, 12'h554, 12'h444, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'haaa, 12'h677, 12'h566, 12'h455, 12'h345, 12'h345, 12'h345, 12'h355, 12'h455, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h445, 12'h345, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h455, 12'h456, 12'h566, 12'h455, 12'h455, 12'h556, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 
12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h456, 12'h455, 12'h456, 12'h677, 12'h899, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hddd, 12'hbbb, 12'h99a, 12'h888, 12'h777, 12'h777, 12'h766, 12'h766, 12'h766, 12'h666, 12'h766, 12'h777, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h667, 12'h677, 12'h778, 12'h888, 12'h99a, 12'hbbb, 12'hccd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbcc, 12'hbbb, 12'haab, 12'haaa, 12'h99a, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h79a, 12'h789, 12'h789, 12'h678, 12'h678, 12'h678, 12'h678, 12'h677, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h788, 12'h788, 12'h788, 12'h788, 12'h788, 12'h788, 
12'h789, 12'h889, 12'h899, 12'h99a, 12'h99a, 12'haaa, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h888, 12'h887, 12'h777, 12'h766, 12'h666, 12'h666, 12'h666, 12'h665, 12'h555, 12'h665, 12'h777, 12'h666, 12'h665, 12'h555, 
12'h554, 12'h554, 12'h555, 12'h665, 12'h666, 12'h665, 12'h655, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h544, 12'h554, 12'h554, 12'h444, 12'h544, 12'h443, 12'h444, 12'h554, 12'h554, 12'h544, 12'h544, 12'h554, 12'h555, 12'h554, 12'h554, 12'h544, 12'h444, 12'h544, 12'h444, 12'h544, 12'h444, 12'h544, 12'h554, 12'h444, 12'h443, 12'h544, 12'h544, 12'h444, 12'h554, 12'h554, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h454, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbcc, 12'h999, 12'h566, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h345, 12'h345, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h355, 12'h355, 12'h455, 12'h455, 12'h355, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h455, 12'h456, 12'h355, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h455, 12'h455, 12'h566, 12'h556, 12'h456, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 
12'h345, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h556, 12'h677, 12'hbbc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h889, 12'h888, 12'h777, 12'h767, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 
12'h665, 12'h666, 12'h666, 12'h665, 12'h655, 12'h665, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h777, 12'h778, 12'h889, 12'haaa, 12'hccc, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hbcc, 12'hbbb, 12'haab, 12'h9aa, 12'h99a, 12'h899, 12'h899, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h79a, 12'h79a, 12'h79a, 12'h78a, 12'h789, 12'h678, 12'h678, 12'h678, 12'h668, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 
12'h778, 12'h778, 12'h788, 12'h889, 12'h889, 12'h99a, 12'h99a, 12'haaa, 12'haab, 12'habb, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hbbb, 12'h888, 12'h887, 12'h777, 12'h776, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h555, 12'h665, 12'h666, 12'h666, 12'h655, 12'h554, 
12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h544, 12'h544, 12'h544, 12'h554, 12'h544, 12'h544, 12'h443, 12'h444, 12'h544, 12'h554, 12'h444, 12'h544, 12'h554, 12'h554, 12'h554, 12'h554, 12'h444, 12'h443, 12'h444, 12'h444, 12'h444, 12'h444, 12'h544, 12'h444, 12'h444, 12'h444, 12'h443, 12'h544, 12'h444, 12'h444, 12'h554, 12'h555, 12'h554, 12'h554, 12'h544, 12'h554, 12'h454, 12'h454, 12'h554, 12'h555, 12'h554, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h788, 12'h999, 12'hbbb, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h455, 12'h345, 12'h345, 12'h245, 12'h234, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h356, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h456, 12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h455, 12'h456, 12'h556, 12'h456, 12'h456, 12'h556, 12'h567, 12'h456, 12'h456, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h455, 12'h455, 12'h455, 12'h345, 12'h445, 12'h455, 12'h455, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h778, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hcdd, 12'hccc, 12'haaa, 12'h878, 12'h878, 12'h888, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h655, 
12'h665, 12'h665, 12'h665, 12'h655, 12'h655, 12'h665, 12'h666, 12'h665, 12'h665, 12'h665, 12'h655, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h667, 12'h777, 12'h888, 12'h999, 12'hbbc, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'h9aa, 12'h89a, 12'h899, 12'h789, 12'h789, 12'h789, 12'h78a, 12'h79a, 12'h79a, 12'h79a, 12'h78a, 12'h68a, 12'h689, 12'h679, 12'h578, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h577, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 
12'h677, 12'h678, 12'h678, 12'h678, 12'h778, 12'h889, 12'h889, 12'h99a, 12'h99a, 12'h9aa, 12'haaa, 12'haab, 12'hbbb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hcdd, 12'h999, 12'h888, 12'h777, 12'h777, 12'h776, 12'h666, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h666, 12'h776, 12'h666, 12'h665, 12'h554, 
12'h554, 12'h555, 12'h665, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h554, 12'h554, 12'h544, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h444, 12'h544, 12'h544, 12'h544, 12'h544, 12'h444, 12'h554, 12'h544, 12'h554, 12'h555, 12'h554, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h443, 12'h443, 12'h444, 12'h554, 12'h544, 12'h444, 12'h544, 12'h443, 12'h444, 12'h444, 12'h444, 12'h444, 12'h554, 12'h554, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h454, 12'h444, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h566, 12'h566, 12'h555, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h899, 12'h566, 12'h455, 12'h344, 12'h345, 12'h245, 12'h345, 12'h345, 12'h345, 12'h355, 12'h345, 12'h346, 12'h456, 12'h456, 12'h356, 12'h456, 12'h456, 12'h457, 12'h457, 12'h456, 12'h456, 12'h457, 12'h567, 12'h467, 12'h457, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h456, 12'h456, 12'h456, 12'h355, 12'h455, 12'h456, 12'h456, 12'h456, 12'h566, 12'h566, 12'h567, 12'h566, 12'h556, 12'h456, 12'h566, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h355, 12'h455, 12'h456, 12'h456, 12'h455, 12'h445, 12'h455, 12'h455, 12'h455, 
12'h455, 12'h455, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h567, 12'h999, 12'hccd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcc, 12'hbbb, 12'hbbb, 12'h999, 12'h767, 12'h777, 12'h777, 12'h776, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h655, 
12'h655, 12'h655, 12'h655, 12'h655, 12'h655, 12'h665, 12'h666, 12'h665, 12'h666, 12'h665, 12'h655, 12'h655, 12'h655, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h777, 12'h777, 12'h778, 12'h999, 12'habb, 12'hccd, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haab, 12'h9aa, 12'h99a, 12'h899, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h78a, 12'h78a, 12'h78a, 12'h68a, 12'h68a, 12'h679, 12'h579, 12'h578, 12'h568, 12'h567, 12'h467, 12'h457, 12'h457, 12'h557, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h467, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h467, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 
12'h567, 12'h667, 12'h667, 12'h668, 12'h678, 12'h778, 12'h789, 12'h889, 12'h889, 12'h899, 12'h99a, 12'h99a, 12'haaa, 12'haab, 12'hbbb, 12'hbcc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'hddd, 12'h999, 12'h777, 12'h777, 12'h877, 12'h776, 12'h666, 12'h665, 12'h665, 12'h665, 12'h555, 12'h554, 12'h555, 12'h776, 12'h777, 12'h666, 12'h665, 12'h555, 
12'h555, 12'h665, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h544, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h544, 12'h554, 12'h554, 12'h444, 12'h554, 12'h544, 12'h554, 12'h554, 12'h555, 12'h555, 12'h554, 12'h544, 12'h444, 12'h554, 12'h544, 12'h444, 12'h444, 12'h444, 12'h544, 12'h544, 12'h444, 12'h444, 12'h443, 12'h443, 12'h443, 12'h444, 12'h443, 12'h444, 12'h443, 12'h443, 12'h443, 12'h443, 12'h443, 12'h544, 12'h554, 12'h454, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h566, 12'h666, 12'h777, 12'h777, 12'h888, 12'haaa, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbcc, 12'h888, 12'h556, 12'h345, 12'h244, 12'h345, 12'h345, 12'h345, 12'h346, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h467, 12'h467, 12'h467, 12'h467, 12'h467, 12'h567, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h568, 12'h567, 12'h568, 12'h567, 12'h467, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h677, 12'h567, 12'h556, 12'h556, 12'h556, 12'h566, 12'h456, 12'h456, 12'h556, 12'h455, 12'h455, 12'h456, 12'h566, 12'h566, 12'h456, 12'h455, 12'h355, 12'h455, 12'h355, 12'h456, 
12'h455, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h455, 12'h455, 12'h445, 12'h345, 12'h355, 12'h456, 12'h556, 12'h778, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hddd, 12'hccc, 12'h99a, 12'h999, 12'h889, 12'h777, 12'h666, 12'h766, 12'h776, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h655, 
12'h655, 12'h555, 12'h655, 12'h655, 12'h655, 12'h665, 12'h666, 12'h666, 12'h666, 12'h665, 12'h655, 12'h555, 12'h555, 12'h655, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h778, 12'h899, 12'h9aa, 12'hbcc, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haab, 12'haaa, 12'haaa, 12'haaa, 12'h9aa, 12'h99a, 12'h99a, 12'h899, 12'h889, 12'h789, 12'h789, 12'h679, 12'h689, 12'h78a, 12'h78a, 12'h78a, 12'h68a, 12'h68a, 12'h67a, 12'h579, 12'h579, 12'h579, 12'h568, 12'h568, 12'h568, 12'h567, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h567, 12'h567, 12'h457, 12'h457, 12'h467, 12'h466, 12'h567, 12'h567, 12'h567, 12'h556, 
12'h557, 12'h567, 12'h567, 12'h567, 12'h667, 12'h668, 12'h778, 12'h778, 12'h789, 12'h889, 12'h889, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'habb, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hded, 12'haba, 12'h777, 12'h777, 12'h776, 12'h887, 12'h776, 12'h666, 12'h666, 12'h655, 12'h665, 12'h665, 12'h555, 12'h655, 12'h666, 12'h776, 12'h665, 12'h665, 12'h655, 
12'h655, 12'h665, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h544, 12'h544, 12'h544, 12'h554, 12'h554, 12'h554, 12'h544, 12'h544, 12'h554, 12'h554, 12'h554, 12'h444, 12'h544, 12'h555, 12'h555, 12'h555, 12'h554, 12'h444, 12'h554, 12'h555, 12'h554, 12'h444, 12'h544, 12'h554, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h443, 12'h444, 12'h444, 12'h443, 12'h444, 12'h443, 12'h443, 12'h443, 12'h444, 12'h444, 12'h444, 12'h555, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h677, 12'h777, 12'h899, 12'habb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'h99a, 12'h667, 12'h455, 12'h244, 12'h234, 12'h245, 12'h345, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h457, 12'h467, 12'h467, 12'h568, 12'h678, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h678, 12'h678, 12'h789, 12'h789, 12'h789, 12'h689, 12'h789, 12'h679, 12'h678, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h456, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h566, 12'h456, 12'h566, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h566, 12'h566, 12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 
12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h455, 12'h456, 12'h456, 12'h566, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h777, 12'h777, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h655, 
12'h555, 12'h655, 12'h655, 12'h655, 12'h655, 12'h665, 12'h665, 12'h666, 12'h666, 12'h666, 12'h665, 12'h655, 12'h555, 12'h655, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h776, 12'h676, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h778, 12'h889, 12'habb, 12'hcdd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'hbbc, 12'haab, 12'h99a, 12'h999, 12'h899, 12'h899, 12'h899, 12'h889, 12'h789, 12'h789, 12'h789, 12'h679, 12'h679, 12'h679, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h67a, 12'h579, 12'h579, 12'h568, 12'h568, 12'h568, 12'h568, 12'h567, 12'h567, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h466, 12'h567, 12'h557, 12'h456, 
12'h456, 12'h457, 12'h557, 12'h557, 12'h567, 12'h567, 12'h667, 12'h668, 12'h668, 12'h778, 12'h678, 12'h678, 12'h788, 12'h789, 12'h899, 12'h99a, 12'haaa, 12'hbbb, 12'hbcc, 12'hccd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h777, 12'h776, 12'h776, 12'h777, 12'h766, 12'h665, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h666, 12'h776, 12'h665, 12'h555, 12'h555, 
12'h665, 12'h665, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h554, 12'h554, 12'h554, 12'h444, 12'h444, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h454, 12'h555, 12'h555, 12'h554, 12'h454, 12'h554, 12'h554, 12'h444, 12'h444, 12'h444, 12'h544, 12'h444, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h443, 12'h443, 12'h444, 12'h444, 12'h444, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h665, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h999, 12'haaa, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h677, 12'h455, 12'h345, 12'h245, 12'h345, 12'h345, 12'h456, 12'h456, 12'h567, 12'h567, 12'h457, 12'h457, 12'h457, 12'h567, 12'h568, 12'h679, 12'h679, 12'h68a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h679, 12'h678, 12'h668, 12'h567, 12'h567, 12'h567, 12'h467, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h567, 12'h566, 12'h566, 12'h556, 12'h566, 12'h456, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h567, 12'h567, 12'h566, 
12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h355, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h788, 12'hbcc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'hbbb, 12'h999, 12'h999, 12'h889, 12'h778, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h555, 
12'h556, 12'h656, 12'h656, 12'h656, 12'h666, 12'h666, 12'h655, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h655, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h677, 12'h888, 12'habb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h99a, 12'h899, 12'h889, 12'h789, 12'h789, 12'h789, 12'h679, 12'h679, 12'h679, 12'h679, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h679, 12'h579, 12'h579, 12'h568, 12'h568, 12'h568, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h456, 12'h557, 12'h557, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h678, 12'h778, 12'h889, 12'h89a, 12'h9aa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h777, 12'h776, 12'h777, 12'h877, 12'h766, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h666, 12'h555, 12'h554, 12'h554, 
12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h554, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h454, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h566, 12'h566, 12'h666, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hdee, 12'habb, 12'h566, 12'h355, 12'h345, 12'h345, 12'h345, 12'h355, 12'h567, 12'h567, 12'h567, 12'h567, 12'h457, 12'h467, 12'h568, 12'h679, 12'h68a, 12'h78a, 12'h79a, 12'h79b, 12'h78a, 12'h78a, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h89b, 12'h78a, 12'h789, 12'h679, 12'h568, 12'h568, 12'h567, 12'h457, 12'h457, 12'h567, 12'h678, 12'h668, 12'h567, 12'h567, 12'h668, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h567, 12'h567, 12'h556, 12'h567, 12'h567, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 
12'h567, 12'h566, 12'h456, 12'h355, 12'h345, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h778, 12'haaa, 12'hccc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbc, 12'h99a, 12'h888, 12'h888, 12'h777, 12'h766, 12'h766, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h655, 12'h555, 
12'h556, 12'h556, 12'h656, 12'h666, 12'h666, 12'h666, 12'h656, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h677, 12'h677, 12'h788, 12'haab, 12'hcdd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'habb, 12'h9aa, 12'h899, 12'h889, 12'h789, 12'h789, 12'h678, 12'h679, 12'h679, 12'h679, 12'h679, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h679, 12'h579, 12'h568, 12'h568, 12'h468, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h557, 12'h557, 12'h557, 12'h557, 12'h457, 12'h456, 12'h356, 12'h356, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h567, 12'h668, 12'h789, 12'h89a, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h777, 12'h777, 12'h776, 12'h887, 12'h887, 12'h777, 12'h766, 12'h665, 12'h555, 12'h555, 12'h554, 12'h555, 12'h665, 12'h666, 12'h665, 12'h555, 12'h554, 12'h554, 
12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h566, 12'h666, 12'h666, 12'h566, 12'h555, 12'h566, 12'h666, 12'h555, 12'h555, 12'h555, 12'h444, 12'h444, 12'h444, 12'h454, 12'h454, 12'h555, 12'h454, 12'h444, 12'h554, 12'h454, 12'h454, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h566, 12'h555, 12'h555, 12'h566, 12'h666, 12'h677, 12'h777, 12'h888, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'h778, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h566, 12'h567, 12'h567, 12'h457, 12'h457, 12'h357, 12'h568, 12'h679, 12'h78a, 12'h79b, 12'h89b, 12'h89c, 12'h8ac, 12'h89b, 12'h89c, 12'h8ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h78a, 12'h679, 12'h678, 12'h678, 12'h578, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h678, 12'h567, 12'h568, 12'h678, 12'h678, 12'h567, 12'h567, 12'h467, 12'h567, 12'h678, 12'h678, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 
12'h567, 12'h567, 12'h566, 12'h456, 12'h455, 12'h355, 12'h455, 12'h456, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h455, 12'h456, 12'h456, 12'h566, 12'h677, 12'haab, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hddd, 12'hbbb, 12'h889, 12'h888, 12'h777, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h666, 12'h666, 12'h666, 12'h667, 
12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h677, 12'h788, 12'haaa, 12'hccd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'hbbc, 12'haab, 12'h99a, 12'h899, 12'h789, 12'h789, 12'h789, 12'h679, 12'h679, 12'h679, 12'h689, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h58a, 12'h58a, 12'h579, 12'h579, 12'h569, 12'h468, 12'h458, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h457, 12'h456, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h456, 12'h456, 12'h557, 12'h456, 12'h557, 12'h557, 12'h557, 12'h457, 12'h567, 12'h678, 12'h789, 12'h899, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h888, 12'h888, 12'h887, 12'h777, 12'h666, 12'h555, 12'h555, 12'h554, 12'h554, 12'h655, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 
12'h555, 12'h555, 12'h565, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h555, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h555, 12'h565, 12'h555, 12'h665, 12'h656, 12'h666, 12'h665, 12'h666, 12'h665, 12'h555, 12'h565, 12'h556, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h666, 12'h666, 12'h666, 12'h677, 12'h888, 12'h999, 12'hbbb, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdd, 12'haaa, 12'h556, 12'h345, 12'h355, 12'h455, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h457, 12'h356, 12'h467, 12'h579, 12'h68a, 12'h79b, 12'h89b, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ad, 12'h9bd, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h79a, 12'h78a, 12'h689, 12'h78a, 12'h679, 12'h679, 12'h578, 12'h578, 12'h678, 12'h679, 12'h789, 12'h789, 12'h789, 12'h679, 12'h678, 12'h678, 12'h679, 12'h678, 12'h568, 12'h568, 12'h568, 12'h678, 12'h678, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 
12'h678, 12'h678, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h355, 12'h455, 12'h456, 12'h556, 12'h567, 12'h788, 12'hbbc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccc, 12'hbcc, 12'hbbb, 12'h99a, 12'h999, 12'h888, 12'h777, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h667, 12'h667, 12'h667, 12'h778, 12'h779, 12'h779, 12'h779, 
12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h767, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h777, 12'h788, 12'haaa, 12'hcdd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h99a, 12'h889, 12'h889, 12'h789, 12'h789, 12'h779, 12'h679, 12'h679, 12'h689, 12'h689, 12'h679, 12'h679, 12'h57a, 12'h58a, 12'h58a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h58a, 12'h57a, 12'h579, 12'h569, 12'h468, 12'h468, 12'h458, 12'h467, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h678, 12'h789, 12'h89a, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'h666, 12'h666, 12'h777, 12'h776, 12'h666, 12'h887, 12'h888, 12'h887, 12'h777, 12'h777, 12'h665, 12'h555, 12'h555, 12'h554, 12'h665, 12'h665, 12'h655, 12'h555, 12'h555, 12'h655, 
12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h666, 12'h665, 12'h665, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h777, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h556, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h777, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h788, 12'h456, 12'h345, 12'h345, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h457, 12'h457, 12'h467, 12'h679, 12'h79b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h79b, 12'h78a, 12'h89b, 12'h89a, 12'h78a, 12'h68a, 12'h689, 12'h68a, 12'h78a, 12'h89a, 12'h89a, 12'h89b, 12'h78a, 12'h789, 12'h78a, 12'h78a, 12'h689, 12'h679, 12'h689, 12'h789, 12'h679, 12'h678, 12'h567, 12'h568, 12'h678, 12'h678, 12'h679, 12'h789, 
12'h789, 12'h789, 12'h678, 12'h567, 12'h467, 12'h457, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h456, 12'h566, 12'h677, 12'hbcc, 12'hdee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'hbbc, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h888, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h668, 12'h779, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 
12'h889, 12'h789, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h767, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h556, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h777, 12'h778, 12'h888, 12'haab, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h9aa, 12'h899, 12'h889, 12'h889, 12'h889, 12'h789, 12'h789, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h579, 12'h579, 12'h579, 12'h57a, 12'h58a, 12'h58a, 12'h68a, 12'h68b, 12'h68b, 12'h68a, 12'h57a, 12'h57a, 12'h579, 12'h579, 12'h569, 12'h468, 12'h468, 12'h457, 12'h457, 12'h457, 12'h457, 12'h356, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h679, 12'h789, 12'h89a, 12'h99a, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h766, 12'h665, 12'h666, 12'h777, 12'h776, 12'h666, 12'h887, 12'h887, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h655, 12'h555, 12'h555, 12'h666, 
12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h667, 12'h777, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h677, 12'h778, 12'h678, 12'h678, 12'h678, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h677, 12'h667, 12'h667, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h566, 12'h566, 12'h566, 12'h556, 12'h565, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h567, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h457, 12'h457, 12'h568, 12'h78a, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h79a, 12'h89b, 12'h79a, 12'h78a, 12'h679, 12'h579, 12'h679, 12'h679, 12'h689, 12'h789, 12'h78a, 
12'h78a, 12'h78a, 12'h689, 12'h678, 12'h578, 12'h567, 12'h456, 12'h456, 12'h355, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h667, 12'h9aa, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h778, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h556, 12'h557, 12'h667, 12'h678, 12'h78a, 12'h88a, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h88a, 12'h78a, 12'h789, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h778, 12'h778, 12'h778, 12'h678, 12'h677, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h777, 12'h778, 12'h788, 12'haab, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccd, 12'hbbb, 12'haaa, 12'h899, 12'h889, 12'h789, 12'h789, 12'h789, 12'h789, 12'h679, 12'h678, 12'h678, 12'h678, 12'h678, 12'h579, 12'h579, 12'h579, 12'h579, 12'h68a, 12'h68a, 12'h68a, 12'h68b, 12'h68b, 12'h68b, 12'h68a, 12'h57a, 12'h57a, 12'h579, 12'h579, 12'h569, 12'h468, 12'h468, 12'h458, 12'h457, 12'h457, 12'h457, 12'h356, 12'h346, 12'h356, 12'h456, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h457, 12'h567, 12'h567, 12'h568, 12'h568, 12'h679, 12'h679, 12'h789, 12'h89a, 12'h9aa, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h887, 12'h666, 12'h665, 12'h665, 12'h776, 12'h777, 12'h776, 12'h777, 12'h777, 12'h777, 12'h776, 12'h777, 12'h777, 12'h777, 12'h766, 12'h666, 12'h665, 12'h655, 12'h655, 12'h666, 12'h666, 12'h666, 
12'h666, 12'h666, 12'h677, 12'h777, 12'h777, 12'h667, 12'h677, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h778, 12'h778, 12'h778, 12'h788, 12'h788, 12'h788, 12'h788, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h788, 12'h789, 12'h788, 12'h788, 12'h778, 12'h778, 12'h789, 12'h778, 12'h778, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h778, 12'h678, 12'h678, 12'h678, 12'h677, 12'h667, 12'h667, 12'h667, 12'h677, 12'h667, 12'h667, 12'h666, 12'h666, 12'h566, 12'h566, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h566, 12'h666, 12'h777, 12'h999, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbc, 12'h788, 12'h556, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h467, 12'h457, 12'h568, 12'h689, 12'h89b, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'h9bd, 12'habd, 12'habe, 12'habe, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'hacd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h8ac, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h68a, 12'h78a, 12'h78a, 12'h78a, 12'h89a, 12'h89b, 
12'h89b, 12'h89a, 12'h78a, 12'h789, 12'h679, 12'h568, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h456, 12'h667, 12'h889, 12'habb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h9aa, 12'h788, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h567, 12'h557, 12'h678, 12'h88a, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 
12'h88b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h779, 12'h778, 12'h778, 12'h778, 12'h678, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h676, 12'h677, 12'h777, 12'h777, 12'h778, 12'haaa, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbc, 12'haab, 12'h99a, 12'h889, 12'h889, 12'h789, 12'h789, 12'h789, 12'h789, 12'h679, 12'h678, 12'h568, 12'h568, 12'h578, 12'h679, 12'h679, 12'h579, 12'h67a, 12'h68a, 12'h68a, 12'h68b, 12'h68b, 12'h68b, 12'h68b, 12'h68a, 12'h58a, 12'h57a, 12'h57a, 12'h579, 12'h569, 12'h469, 12'h468, 12'h568, 12'h458, 12'h458, 12'h457, 12'h457, 12'h457, 12'h357, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h356, 12'h456, 12'h446, 12'h346, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h556, 12'h557, 12'h557, 12'h557, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h568, 12'h568, 12'h568, 12'h678, 12'h679, 12'h789, 12'h89a, 12'h9aa, 12'haab, 12'hbbb, 12'hccc, 12'hddd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h777, 12'h666, 12'h555, 12'h665, 12'h776, 12'h777, 12'h777, 12'h776, 12'h777, 12'h776, 12'h666, 12'h776, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h655, 12'h655, 12'h666, 12'h666, 12'h666, 
12'h777, 12'h778, 12'h778, 12'h788, 12'h778, 12'h778, 12'h778, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h88a, 12'h789, 12'h789, 12'h789, 12'h79a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h778, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h779, 12'h678, 12'h678, 12'h677, 12'h667, 12'h678, 12'h678, 12'h678, 12'h678, 12'h677, 12'h667, 12'h666, 12'h566, 12'h566, 12'h666, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hddd, 12'heef, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h99a, 12'h677, 12'h556, 12'h456, 12'h455, 12'h456, 12'h456, 12'h456, 12'h567, 12'h467, 12'h457, 12'h567, 12'h679, 12'h79a, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'habe, 12'hace, 12'hace, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hacd, 12'habd, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h79b, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h679, 12'h679, 12'h567, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h355, 12'h345, 12'h345, 12'h456, 12'h456, 12'h667, 12'h889, 12'hbcc, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hccc, 12'habb, 12'h999, 12'h777, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h667, 12'h556, 12'h667, 12'h679, 12'h88a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 
12'h88b, 12'h78b, 12'h78b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h779, 12'h779, 12'h778, 12'h678, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h777, 12'h778, 12'haab, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'habb, 12'h9aa, 12'h89a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h779, 12'h679, 12'h679, 12'h678, 12'h568, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h57a, 12'h68a, 12'h68a, 12'h68b, 12'h78b, 12'h79b, 12'h68b, 12'h68b, 12'h58a, 12'h57a, 12'h57a, 12'h479, 12'h469, 12'h469, 12'h468, 12'h468, 12'h458, 12'h468, 12'h458, 12'h458, 12'h457, 12'h458, 12'h458, 12'h458, 12'h457, 12'h457, 12'h457, 12'h357, 12'h356, 12'h356, 12'h356, 12'h356, 12'h456, 12'h456, 12'h346, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h556, 12'h557, 12'h557, 12'h557, 12'h557, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h679, 12'h789, 12'h89a, 12'h99a, 12'h9aa, 12'habb, 12'hbcc, 12'hccd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'haa9, 12'h887, 12'h776, 12'h666, 12'h555, 12'h655, 12'h777, 12'h777, 12'h777, 12'h776, 12'h776, 12'h666, 12'h666, 12'h666, 12'h766, 12'h776, 12'h776, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 
12'h777, 12'h778, 12'h788, 12'h788, 12'h788, 12'h789, 12'h789, 12'h78a, 12'h78a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h79a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89a, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h78a, 12'h79a, 12'h79a, 12'h79a, 12'h79a, 12'h78a, 12'h79a, 12'h79a, 12'h79b, 12'h89b, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h779, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h678, 12'h678, 12'h666, 12'h566, 12'h566, 12'h566, 12'h556, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h566, 12'h566, 12'h555, 12'h555, 12'h555, 12'h444, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'h999, 12'hbbb, 12'heee, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h677, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h466, 12'h567, 12'h567, 12'h567, 12'h568, 12'h689, 12'h89b, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'habe, 12'hace, 12'hace, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h89b, 12'h89c, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h568, 12'h467, 12'h456, 12'h456, 12'h456, 12'h355, 12'h355, 12'h355, 12'h345, 12'h455, 12'h456, 12'h566, 12'h778, 12'h9aa, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcc, 12'haaa, 12'h999, 12'h888, 12'h787, 12'h777, 12'h666, 12'h666, 12'h567, 12'h667, 12'h668, 12'h88a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 
12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h78b, 12'h78b, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h779, 12'h778, 12'h778, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h776, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h565, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h778, 12'h889, 12'hbbb, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccd, 12'hbbc, 12'haab, 12'h99a, 12'h889, 12'h789, 12'h789, 12'h779, 12'h679, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h57a, 12'h68a, 12'h68b, 12'h68b, 12'h79b, 12'h69b, 12'h68b, 12'h68b, 12'h58a, 12'h68a, 12'h67a, 12'h57a, 12'h469, 12'h469, 12'h469, 12'h468, 12'h468, 12'h468, 12'h468, 12'h468, 12'h568, 12'h568, 12'h568, 12'h468, 12'h568, 12'h468, 12'h457, 12'h357, 12'h357, 12'h357, 12'h356, 12'h356, 12'h356, 12'h456, 12'h346, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h457, 12'h567, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h789, 12'h89a, 12'h89a, 12'h99a, 12'haab, 12'hbbc, 12'hcdd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h777, 12'h666, 12'h665, 12'h555, 12'h665, 12'h777, 12'h777, 12'h877, 12'h777, 12'h666, 12'h666, 12'h666, 12'h776, 12'h666, 12'h766, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 
12'h778, 12'h778, 12'h788, 12'h789, 12'h789, 12'h789, 12'h78a, 12'h79a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79a, 12'h79a, 12'h79a, 12'h79a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h678, 12'h678, 12'h779, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h677, 12'h566, 12'h666, 12'h555, 12'h566, 12'h566, 12'h566, 12'h555, 12'h555, 12'h455, 12'h444, 12'h455, 12'h455, 12'h555, 12'h555, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'haaa, 12'hddd, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h567, 12'h556, 12'h456, 12'h355, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h467, 12'h567, 12'h678, 12'h79a, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h89c, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 
12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89b, 12'h79b, 12'h78a, 12'h679, 12'h568, 12'h457, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h345, 12'h456, 12'h556, 12'h667, 12'h899, 12'hcdd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'habb, 12'h889, 12'h777, 12'h777, 12'h677, 12'h667, 12'h666, 12'h566, 12'h667, 12'h789, 12'h99b, 12'h9ac, 12'haac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h8ac, 
12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h78b, 12'h78b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h78a, 12'h789, 12'h778, 12'h678, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h565, 12'h565, 12'h666, 12'h666, 12'h666, 12'h776, 12'h666, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h777, 12'h778, 12'h99a, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcc, 12'habb, 12'h9aa, 12'h89a, 12'h789, 12'h789, 12'h679, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h679, 12'h679, 12'h579, 12'h679, 12'h68a, 12'h68a, 12'h68b, 12'h68b, 12'h79b, 12'h78b, 12'h68b, 12'h68b, 12'h68a, 12'h68a, 12'h68a, 12'h57a, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h679, 12'h679, 12'h679, 12'h679, 12'h579, 12'h569, 12'h568, 12'h568, 12'h457, 12'h457, 12'h457, 12'h357, 12'h456, 12'h356, 12'h456, 12'h456, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h457, 12'h567, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h789, 12'h889, 12'h899, 12'h99a, 12'haab, 12'hbcc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h776, 12'h666, 12'h665, 12'h555, 12'h665, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h766, 12'h777, 12'h777, 12'h778, 12'h888, 12'h889, 12'h889, 12'h889, 12'h788, 12'h778, 
12'h788, 12'h789, 12'h789, 12'h889, 12'h789, 12'h78a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h679, 12'h779, 12'h689, 12'h679, 12'h679, 12'h679, 12'h689, 12'h789, 12'h778, 12'h566, 12'h556, 12'h566, 12'h555, 12'h556, 12'h667, 12'h565, 12'h555, 12'h555, 12'h455, 12'h444, 12'h444, 12'h455, 12'h555, 12'h566, 12'h555, 12'h455, 12'h555, 12'h454, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h999, 12'hccc, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'h567, 12'h556, 12'h345, 12'h345, 12'h456, 12'h456, 12'h567, 12'h567, 12'h467, 12'h467, 12'h568, 12'h78a, 12'h8ab, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h9bd, 12'habd, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habe, 12'hbce, 12'hace, 12'habd, 12'habd, 12'hace, 12'habe, 12'habe, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 
12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h79b, 12'h78a, 12'h679, 12'h568, 12'h467, 12'h456, 12'h456, 12'h456, 12'h455, 12'h345, 12'h355, 12'h456, 12'h456, 12'h567, 12'h788, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcc, 12'haaa, 12'h889, 12'h677, 12'h667, 12'h667, 12'h667, 12'h567, 12'h668, 12'h88a, 12'h9ac, 12'haac, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 
12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h789, 12'h779, 12'h778, 12'h768, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h565, 12'h665, 12'h665, 12'h666, 12'h666, 12'h777, 12'h777, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h778, 12'h889, 12'hbbb, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h9ab, 12'h89a, 12'h89a, 12'h789, 12'h679, 12'h678, 12'h578, 12'h568, 12'h668, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h68a, 12'h68a, 12'h68a, 12'h68b, 12'h68b, 12'h79b, 12'h79b, 12'h79b, 12'h68b, 12'h68b, 12'h68a, 12'h78a, 12'h68a, 12'h579, 12'h579, 12'h579, 12'h579, 12'h679, 12'h67a, 12'h78a, 12'h79a, 12'h79a, 12'h78a, 12'h679, 12'h679, 12'h579, 12'h568, 12'h468, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h789, 12'h789, 12'h889, 12'h99a, 12'habb, 12'hccc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h777, 12'h776, 12'h666, 12'h665, 12'h655, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h666, 12'h766, 12'h776, 12'h777, 12'h777, 12'h888, 12'h89a, 12'h9ab, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h789, 
12'h889, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h689, 12'h679, 12'h789, 12'h789, 12'h789, 12'h667, 12'h555, 12'h666, 12'h555, 12'h566, 12'h677, 12'h666, 12'h667, 12'h667, 12'h555, 12'h455, 12'h444, 12'h444, 12'h555, 12'h566, 12'h566, 12'h555, 12'h455, 12'h555, 12'h454, 12'h455, 12'h555, 12'h555, 12'h555, 12'h666, 12'h888, 12'hccc, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbcc, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h567, 12'h667, 12'h567, 12'h467, 12'h567, 12'h678, 12'h79a, 12'h8ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h79c, 12'h89c, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'hace, 12'habe, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 
12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h79a, 12'h78a, 12'h679, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h456, 12'h456, 12'h566, 12'h788, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h889, 12'h777, 12'h667, 12'h667, 12'h667, 12'h779, 12'h99b, 12'haac, 12'haac, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h779, 12'h778, 12'h768, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h565, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h677, 12'h778, 12'h99a, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccd, 12'hbbc, 12'haab, 12'h89a, 12'h89a, 12'h789, 12'h789, 12'h678, 12'h578, 12'h568, 12'h568, 12'h568, 12'h678, 12'h668, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h68a, 12'h68a, 12'h68a, 12'h68a, 12'h78a, 12'h79b, 12'h79b, 12'h79b, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h679, 12'h579, 12'h579, 12'h679, 12'h679, 12'h78a, 12'h78a, 12'h89b, 12'h89a, 12'h78a, 12'h68a, 12'h679, 12'h578, 12'h568, 12'h468, 12'h567, 12'h457, 12'h457, 12'h457, 12'h346, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h346, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h468, 12'h568, 12'h568, 12'h568, 12'h567, 12'h568, 12'h678, 12'h779, 12'h789, 12'h899, 12'haaa, 12'hbbc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h776, 12'h666, 12'h777, 12'h777, 12'h888, 12'h889, 12'h89a, 12'h9ab, 12'habc, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 
12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h8ac, 12'h9ab, 12'h9ab, 12'h8ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h89b, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79a, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h689, 12'h789, 12'h789, 12'h789, 12'h677, 12'h555, 12'h566, 12'h555, 12'h667, 12'h778, 12'h678, 12'h789, 12'h678, 12'h666, 12'h555, 12'h444, 12'h444, 12'h444, 12'h555, 12'h565, 12'h555, 12'h454, 12'h555, 12'h454, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h888, 12'hbbb, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h567, 12'h556, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h679, 12'h89b, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9bd, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h78a, 12'h789, 12'h578, 12'h467, 12'h456, 12'h456, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h566, 12'h778, 12'hbcc, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccc, 12'h9aa, 12'h889, 12'h778, 12'h777, 12'h667, 12'h567, 12'h779, 12'h9ab, 12'habc, 12'habc, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h779, 12'h778, 12'h767, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h555, 12'h555, 12'h566, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h666, 12'h666, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h889, 12'haab, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcc, 12'haab, 12'h9aa, 12'h89a, 12'h789, 12'h789, 12'h679, 12'h678, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h668, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h689, 12'h689, 12'h689, 12'h689, 12'h68a, 12'h68a, 12'h78a, 12'h78a, 12'h78a, 12'h68a, 12'h689, 12'h679, 12'h679, 12'h679, 12'h569, 12'h579, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h689, 12'h679, 12'h579, 12'h568, 12'h568, 12'h468, 12'h457, 12'h457, 12'h457, 12'h457, 12'h347, 12'h446, 12'h446, 12'h446, 12'h446, 12'h346, 12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h346, 12'h346, 12'h346, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h568, 12'h567, 12'h568, 12'h568, 12'h678, 12'h678, 12'h789, 12'h99a, 12'habb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h666, 12'h665, 12'h666, 12'h776, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h776, 12'h777, 12'h888, 12'h889, 12'h89a, 12'h9ab, 12'habc, 12'habd, 12'habc, 12'h9ab, 12'habc, 12'hbcd, 12'habd, 
12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79a, 12'h79b, 12'h79b, 12'h79b, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h78a, 12'h789, 12'h689, 12'h677, 12'h556, 12'h567, 12'h678, 12'h789, 12'h78a, 12'h79a, 12'h79a, 12'h789, 12'h678, 12'h666, 12'h555, 12'h455, 12'h444, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h454, 12'h455, 12'h555, 12'h555, 12'h555, 12'h666, 12'h888, 12'hbbb, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h889, 12'h567, 12'h456, 12'h456, 12'h456, 12'h566, 12'h567, 12'h456, 12'h567, 12'h567, 12'h678, 12'h78a, 12'h89b, 12'h9ac, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'habe, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'hace, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h78a, 12'h679, 12'h567, 12'h456, 12'h456, 12'h456, 12'h455, 12'h355, 12'h455, 12'h456, 12'h556, 12'h788, 12'hccc, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h778, 12'h677, 12'h667, 12'h667, 12'h789, 12'h9ab, 12'habc, 12'habc, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habd, 12'habe, 12'habd, 12'habd, 
12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h779, 12'h778, 12'h778, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h666, 12'h555, 12'h555, 12'h556, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h778, 12'h99a, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'habb, 12'h9ab, 12'h89a, 12'h789, 12'h689, 12'h689, 12'h679, 12'h678, 12'h568, 12'h567, 12'h567, 12'h567, 12'h568, 12'h668, 12'h678, 12'h678, 12'h779, 12'h779, 12'h779, 12'h789, 12'h789, 12'h679, 12'h679, 12'h679, 12'h689, 12'h689, 12'h679, 12'h679, 12'h679, 12'h678, 12'h679, 12'h678, 12'h668, 12'h668, 12'h568, 12'h568, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h68a, 12'h679, 12'h579, 12'h569, 12'h568, 12'h568, 12'h568, 12'h568, 12'h458, 12'h358, 12'h458, 12'h357, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 
12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h346, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h778, 12'h889, 12'h9aa, 12'hbcc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h665, 12'h665, 12'h666, 12'h776, 12'h776, 12'h776, 12'h777, 12'h777, 12'h877, 12'h777, 12'h766, 12'h776, 12'h777, 12'h888, 12'h778, 12'h899, 12'h9ab, 12'habd, 12'hbcd, 12'hbbd, 12'habc, 12'habc, 12'hbcd, 12'hbcd, 12'habd, 
12'habc, 12'habc, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h689, 12'h689, 12'h689, 12'h79a, 12'h8ab, 12'h8ab, 12'h8ab, 12'h8ab, 12'h89b, 12'h79a, 12'h789, 12'h677, 12'h566, 12'h555, 12'h555, 12'h444, 12'h444, 12'h555, 12'h555, 12'h455, 12'h555, 12'h454, 12'h455, 12'h555, 12'h555, 12'h666, 12'h888, 12'hbbb, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h677, 12'h566, 12'h566, 12'h566, 12'h566, 12'h456, 12'h567, 12'h466, 12'h567, 12'h567, 12'h678, 12'h78a, 12'h89b, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habe, 12'hace, 12'hace, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hbdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'habe, 12'habe, 12'hace, 12'habe, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89a, 12'h78a, 12'h678, 12'h567, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h456, 12'h556, 12'h778, 12'hbbc, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h677, 12'h567, 12'h567, 12'h789, 12'h9ab, 12'haac, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h789, 12'h779, 12'h778, 12'h778, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h889, 12'haab, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'hbbc, 12'haab, 12'h99a, 12'h78a, 12'h689, 12'h679, 12'h679, 12'h678, 12'h578, 12'h567, 12'h567, 12'h567, 12'h567, 12'h668, 12'h678, 12'h678, 12'h778, 12'h789, 12'h789, 12'h789, 12'h778, 12'h678, 12'h568, 12'h568, 12'h678, 12'h678, 12'h678, 12'h567, 12'h467, 12'h467, 12'h567, 12'h568, 12'h568, 12'h568, 12'h668, 12'h679, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h689, 12'h579, 12'h568, 12'h468, 12'h568, 12'h568, 12'h579, 12'h579, 12'h569, 12'h568, 12'h568, 12'h568, 12'h568, 12'h558, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 
12'h446, 12'h446, 12'h346, 12'h346, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h346, 12'h446, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h567, 12'h568, 12'h678, 12'h789, 12'h99a, 12'hbbb, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h888, 12'h666, 12'h665, 12'h665, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h887, 12'h766, 12'h777, 12'h778, 12'h888, 12'h889, 12'h9aa, 12'habc, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'hbce, 12'hbcd, 12'hbcd, 12'hbcd, 
12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h78a, 12'h78a, 12'h78a, 12'h79b, 12'h8ab, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h89b, 12'h79a, 12'h789, 12'h677, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h454, 12'h444, 12'h555, 12'h555, 12'h555, 12'h666, 12'h788, 12'habb, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h679, 12'h89a, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'habd, 12'habe, 12'hace, 12'hace, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hbdf, 12'hbdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'habe, 12'hace, 12'habe, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h79a, 12'h678, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h788, 12'hbbc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hbbb, 12'h889, 12'h778, 12'h667, 12'h557, 12'h779, 12'h9ab, 12'habc, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h88b, 12'h88a, 12'h779, 12'h779, 12'h778, 12'h777, 12'h767, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h766, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbbc, 12'habb, 12'h9ab, 12'h89a, 12'h789, 12'h689, 12'h679, 12'h678, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h668, 12'h678, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h668, 12'h567, 12'h457, 12'h466, 12'h567, 12'h567, 12'h567, 12'h457, 12'h457, 12'h457, 12'h557, 12'h668, 12'h678, 12'h679, 12'h779, 12'h789, 12'h78a, 12'h78a, 12'h78a, 12'h68a, 12'h579, 12'h569, 12'h468, 12'h468, 12'h468, 12'h568, 12'h679, 12'h68a, 12'h679, 12'h679, 12'h679, 12'h679, 12'h569, 12'h568, 12'h568, 12'h567, 12'h457, 12'h567, 12'h567, 12'h567, 12'h557, 12'h557, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 
12'h446, 12'h446, 12'h346, 12'h345, 12'h346, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h446, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h468, 12'h568, 12'h568, 12'h568, 12'h568, 12'h467, 12'h567, 12'h567, 12'h678, 12'h788, 12'h899, 12'haab, 12'hccc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h777, 12'h666, 12'h666, 12'h666, 12'h776, 12'h777, 12'h777, 12'h877, 12'h877, 12'h887, 12'h888, 12'h777, 12'h777, 12'h777, 12'h788, 12'h889, 12'h9aa, 12'habc, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hacd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h89b, 12'h79a, 12'h688, 12'h667, 12'h566, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h454, 12'h444, 12'h455, 12'h555, 12'h555, 12'h566, 12'h777, 12'haaa, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h677, 12'h556, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h689, 12'h89b, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hbde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'h9bd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h89b, 12'h679, 12'h567, 12'h467, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h788, 12'hccc, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haab, 12'h788, 12'h667, 12'h667, 12'h779, 12'h9ab, 12'habc, 12'habc, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h779, 12'h778, 12'h778, 12'h777, 12'h767, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h999, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcc, 12'habb, 12'h9ab, 12'h89a, 12'h789, 12'h679, 12'h678, 12'h678, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h668, 12'h678, 12'h678, 12'h678, 12'h668, 12'h667, 12'h567, 12'h557, 12'h456, 12'h456, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h557, 12'h557, 12'h568, 12'h678, 12'h779, 12'h78a, 12'h78a, 12'h78a, 12'h689, 12'h679, 12'h679, 12'h679, 12'h569, 12'h468, 12'h468, 12'h568, 12'h579, 12'h679, 12'h68a, 12'h78a, 12'h68a, 12'h679, 12'h679, 12'h679, 12'h679, 12'h579, 12'h668, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h678, 12'h668, 12'h567, 12'h456, 12'h456, 12'h446, 12'h446, 
12'h446, 12'h446, 12'h346, 12'h346, 12'h446, 12'h446, 12'h445, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h446, 12'h456, 12'h457, 12'h457, 12'h357, 12'h357, 12'h468, 12'h568, 12'h568, 12'h568, 12'h568, 12'h457, 12'h457, 12'h567, 12'h567, 12'h678, 12'h889, 12'h9aa, 12'hbbc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h887, 12'h766, 12'h666, 12'h666, 12'h666, 12'h776, 12'h777, 12'h777, 12'h887, 12'h888, 12'h887, 12'h888, 12'h777, 12'h777, 12'h778, 12'h888, 12'h89a, 12'habc, 12'hbcd, 12'hbcd, 12'hbce, 12'hbcd, 12'habd, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h7ac, 12'h7ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h79a, 12'h789, 12'h678, 12'h666, 12'h666, 12'h555, 12'h455, 12'h555, 12'h555, 12'h455, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h777, 12'haaa, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h778, 12'h566, 12'h566, 12'h456, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h78a, 12'h8ab, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 
12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h89b, 12'h789, 12'h578, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h678, 12'hbcc, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdee, 12'hbbc, 12'h99a, 12'h778, 12'h668, 12'h789, 12'h9ab, 12'habc, 12'habd, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h88a, 12'h779, 12'h779, 12'h778, 12'h778, 12'h777, 12'h767, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h888, 12'haab, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'habb, 12'haaa, 12'h89a, 12'h789, 12'h789, 12'h678, 12'h578, 12'h578, 12'h568, 12'h567, 12'h457, 12'h557, 12'h557, 12'h557, 12'h567, 12'h667, 12'h567, 12'h567, 12'h557, 12'h557, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h556, 12'h456, 12'h556, 12'h557, 12'h668, 12'h779, 12'h789, 12'h789, 12'h789, 12'h679, 12'h679, 12'h568, 12'h568, 12'h579, 12'h679, 12'h579, 12'h579, 12'h579, 12'h679, 12'h679, 12'h68a, 12'h68a, 12'h679, 12'h579, 12'h579, 12'h679, 12'h579, 12'h579, 12'h568, 12'h568, 12'h567, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h668, 12'h567, 12'h556, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h467, 12'h457, 12'h567, 12'h567, 12'h678, 12'h788, 12'h99a, 12'hbbb, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h999, 12'h777, 12'h666, 12'h766, 12'h766, 12'h766, 12'h777, 12'h877, 12'h777, 12'h888, 12'h888, 12'h887, 12'h888, 12'h777, 12'h777, 12'h778, 12'h889, 12'h9ab, 12'hbcd, 12'hbce, 12'hbce, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hbce, 12'hbce, 12'hace, 12'hacd, 12'hacd, 12'habd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h7ac, 12'h7ac, 12'h7ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8bc, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h89b, 12'h78a, 12'h788, 12'h666, 12'h666, 12'h566, 12'h455, 12'h555, 12'h555, 12'h555, 12'h445, 12'h555, 12'h555, 12'h555, 12'h555, 12'h777, 12'haaa, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h778, 12'h556, 12'h556, 12'h566, 12'h567, 12'h456, 12'h566, 12'h567, 12'h678, 12'h679, 12'h89a, 12'h9ac, 12'h9bc, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 
12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h789, 12'h678, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h9aa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'haab, 12'h788, 12'h668, 12'h679, 12'h99b, 12'haac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h99c, 12'h89b, 12'h88a, 12'h78a, 12'h779, 12'h779, 12'h778, 12'h778, 12'h777, 12'h767, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h999, 12'hbbc, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbbb, 12'haaa, 12'h99a, 12'h889, 12'h789, 12'h678, 12'h678, 12'h568, 12'h568, 12'h567, 12'h457, 12'h457, 12'h556, 12'h556, 12'h556, 12'h557, 12'h557, 12'h557, 12'h557, 12'h557, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h556, 12'h557, 12'h557, 12'h667, 12'h778, 12'h779, 12'h779, 12'h678, 12'h668, 12'h568, 12'h568, 12'h468, 12'h568, 12'h579, 12'h679, 12'h579, 12'h579, 12'h579, 12'h679, 12'h679, 12'h679, 12'h579, 12'h579, 12'h579, 12'h569, 12'h569, 12'h569, 12'h568, 12'h568, 12'h457, 12'h457, 12'h457, 12'h456, 12'h567, 12'h667, 12'h668, 12'h567, 12'h557, 12'h556, 12'h456, 12'h456, 
12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h446, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h568, 12'h568, 12'h457, 12'h457, 12'h567, 12'h567, 12'h678, 12'h788, 12'h999, 12'habb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h887, 12'h887, 12'h888, 12'h787, 12'h777, 12'h888, 12'h777, 12'h777, 12'h788, 12'h89a, 12'habc, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcde, 12'hbce, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8bc, 12'h8bc, 12'h9bc, 12'h8ac, 12'h8ac, 12'h89b, 12'h79a, 12'h789, 12'h677, 12'h666, 12'h666, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h455, 12'h555, 12'h555, 12'h555, 12'h677, 12'haaa, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h778, 12'h556, 12'h566, 12'h567, 12'h566, 12'h566, 12'h466, 12'h567, 12'h678, 12'h779, 12'h89b, 12'h9ac, 12'h9bc, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 
12'h9bd, 12'h9bd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h78a, 12'h678, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h9aa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h99a, 12'h678, 12'h678, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h99c, 12'h89b, 12'h88a, 12'h78a, 12'h779, 12'h778, 12'h778, 12'h778, 12'h777, 12'h767, 12'h667, 12'h667, 12'h667, 12'h666, 12'h677, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbc, 12'haab, 12'h99a, 12'h889, 12'h789, 12'h678, 12'h678, 12'h568, 12'h568, 12'h567, 12'h567, 12'h457, 12'h456, 12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h457, 12'h556, 12'h557, 12'h557, 12'h567, 12'h667, 12'h678, 12'h778, 12'h678, 12'h678, 12'h568, 12'h567, 12'h568, 12'h468, 12'h468, 12'h568, 12'h579, 12'h579, 12'h569, 12'h569, 12'h569, 12'h679, 12'h679, 12'h579, 12'h579, 12'h579, 12'h579, 12'h569, 12'h569, 12'h568, 12'h568, 12'h457, 12'h357, 12'h346, 12'h346, 12'h346, 12'h346, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 
12'h456, 12'h557, 12'h557, 12'h557, 12'h556, 12'h456, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h446, 12'h456, 12'h456, 12'h457, 12'h457, 12'h457, 12'h557, 12'h568, 12'h568, 12'h568, 12'h568, 12'h467, 12'h457, 12'h457, 12'h567, 12'h567, 12'h678, 12'h778, 12'h899, 12'haaa, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h777, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h887, 12'h777, 12'h777, 12'h787, 12'h777, 12'h877, 12'h777, 12'h788, 12'h889, 12'h9ab, 12'hbcd, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hbce, 12'hbde, 12'hbde, 12'hbde, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9bc, 12'h9bc, 12'h8bc, 12'h8bc, 12'h8ac, 12'h8ab, 12'h89a, 12'h789, 12'h677, 12'h666, 12'h566, 12'h565, 12'h455, 12'h555, 12'h565, 12'h555, 12'h555, 12'h555, 12'h565, 12'h555, 12'h677, 12'h9aa, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'h899, 12'h567, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h789, 12'h89b, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hace, 12'hacd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habe, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 
12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h79a, 12'h689, 12'h577, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdee, 12'habb, 12'h788, 12'h678, 12'h88a, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h99c, 12'h89b, 12'h88b, 12'h88a, 12'h789, 12'h779, 12'h778, 12'h778, 12'h778, 12'h777, 12'h767, 12'h777, 12'h677, 12'h667, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h999, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccc, 12'habb, 12'h99a, 12'h889, 12'h789, 12'h778, 12'h678, 12'h668, 12'h568, 12'h568, 12'h567, 12'h557, 12'h456, 12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h557, 12'h667, 12'h667, 12'h667, 12'h567, 12'h557, 12'h557, 12'h457, 12'h457, 12'h557, 12'h567, 12'h667, 12'h668, 12'h678, 12'h678, 12'h678, 12'h668, 12'h568, 12'h568, 12'h568, 12'h468, 12'h468, 12'h568, 12'h579, 12'h579, 12'h579, 12'h469, 12'h469, 12'h569, 12'h579, 12'h679, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h569, 12'h568, 12'h568, 12'h457, 12'h457, 12'h456, 12'h346, 12'h346, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h446, 
12'h456, 12'h556, 12'h557, 12'h557, 12'h557, 12'h456, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h445, 12'h446, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h568, 12'h568, 12'h567, 12'h457, 12'h457, 12'h457, 12'h567, 12'h567, 12'h678, 12'h778, 12'h889, 12'h9aa, 12'hbcc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbba, 12'h888, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h878, 12'h777, 12'h777, 12'h877, 12'h888, 12'h89a, 12'habc, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8ac, 12'h8ab, 12'h89b, 12'h79a, 12'h778, 12'h666, 12'h566, 12'h566, 12'h555, 12'h555, 12'h566, 12'h555, 12'h555, 12'h555, 12'h565, 12'h565, 12'h666, 12'h9aa, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'h9aa, 12'h567, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h89a, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'habe, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h89a, 12'h689, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'habb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'h99a, 12'h668, 12'h789, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h99c, 12'h89b, 12'h88a, 12'h78a, 12'h789, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'haaa, 12'h999, 12'h789, 12'h778, 12'h668, 12'h668, 12'h668, 12'h668, 12'h568, 12'h557, 12'h457, 12'h456, 12'h446, 12'h446, 12'h456, 12'h456, 12'h457, 12'h457, 12'h557, 12'h567, 12'h667, 12'h667, 12'h667, 12'h567, 12'h567, 12'h557, 12'h557, 12'h557, 12'h567, 12'h667, 12'h667, 12'h678, 12'h678, 12'h678, 12'h668, 12'h678, 12'h678, 12'h568, 12'h568, 12'h578, 12'h579, 12'h579, 12'h679, 12'h579, 12'h579, 12'h569, 12'h569, 12'h569, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h569, 12'h569, 12'h568, 12'h458, 12'h457, 12'h356, 12'h456, 12'h346, 12'h446, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 
12'h345, 12'h456, 12'h456, 12'h557, 12'h557, 12'h556, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h446, 12'h456, 12'h457, 12'h557, 12'h567, 12'h567, 12'h568, 12'h567, 12'h567, 12'h457, 12'h457, 12'h457, 12'h567, 12'h567, 12'h678, 12'h678, 12'h788, 12'h99a, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h877, 12'h666, 12'h666, 12'h666, 12'h776, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h777, 12'h777, 12'h888, 12'h899, 12'h9ab, 12'habc, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 
12'hcce, 12'hbde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hbce, 12'hace, 12'habd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8bc, 12'h9bd, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8ac, 12'h8ac, 12'h89b, 12'h79a, 12'h789, 12'h667, 12'h555, 12'h566, 12'h566, 12'h555, 12'h566, 12'h566, 12'h566, 12'h565, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haab, 12'h567, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h578, 12'h679, 12'h89b, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'hbbd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habd, 12'habd, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h89a, 12'h789, 12'h567, 12'h566, 12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h567, 12'hbbc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h889, 12'h778, 12'h99b, 12'haac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'hace, 12'hace, 12'hace, 12'hbce, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h89b, 12'h89b, 12'h88a, 12'h789, 12'h789, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h666, 12'h666, 12'h566, 12'h655, 12'h666, 12'h777, 12'h889, 12'haab, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'habb, 12'h99a, 12'h889, 12'h778, 12'h668, 12'h668, 12'h678, 12'h668, 12'h668, 12'h567, 12'h457, 12'h456, 12'h456, 12'h446, 12'h446, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h668, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h667, 12'h678, 12'h778, 12'h778, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h579, 12'h579, 12'h569, 12'h579, 12'h579, 12'h579, 12'h679, 12'h579, 12'h578, 12'h568, 12'h568, 12'h569, 12'h579, 12'h569, 12'h568, 12'h568, 12'h557, 12'h457, 12'h457, 12'h446, 12'h346, 12'h346, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h335, 
12'h345, 12'h446, 12'h456, 12'h556, 12'h456, 12'h456, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h457, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h457, 12'h457, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h788, 12'h999, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h776, 12'h777, 12'h777, 12'h777, 12'h888, 12'h787, 12'h787, 12'h777, 12'h888, 12'h899, 12'h9ab, 12'habc, 12'hbcd, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hbde, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9bd, 12'h9bc, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8bc, 12'h8ac, 12'h8ab, 12'h79a, 12'h789, 12'h677, 12'h566, 12'h556, 12'h566, 12'h565, 12'h565, 12'h566, 12'h666, 12'h566, 12'h565, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haab, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h789, 12'h89b, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h89b, 12'h89a, 12'h89a, 12'h78a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h9ab, 12'habc, 12'habd, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'habd, 12'habd, 12'h9bc, 12'h9ac, 12'h9ac, 12'h8ab, 12'h89a, 12'h789, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'hbcc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'habb, 12'h889, 12'h99a, 12'haab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h78a, 12'h789, 12'h789, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h566, 12'h666, 12'h778, 12'h9aa, 12'hbcc, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbc, 12'haaa, 12'h999, 12'h889, 12'h678, 12'h668, 12'h668, 12'h678, 12'h668, 12'h567, 12'h557, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h678, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h679, 12'h679, 12'h579, 12'h468, 12'h468, 12'h468, 12'h568, 12'h578, 12'h679, 12'h669, 12'h668, 12'h568, 12'h568, 12'h568, 12'h457, 12'h446, 12'h456, 12'h456, 12'h446, 12'h345, 12'h345, 12'h345, 12'h335, 
12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h456, 12'h456, 12'h457, 12'h457, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h778, 12'h889, 12'haab, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h787, 12'h787, 12'h888, 12'h887, 12'h888, 12'h899, 12'h9ab, 12'habc, 12'hbcd, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 
12'hcde, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h8ab, 12'h8ac, 12'h8ac, 12'h8bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h8bc, 12'h9bd, 12'h8bc, 12'h8ac, 12'h8ab, 12'h79a, 12'h689, 12'h677, 12'h677, 12'h566, 12'h566, 12'h566, 12'h565, 12'h566, 12'h566, 12'h566, 12'h565, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h9aa, 12'h567, 12'h567, 12'h567, 12'h677, 12'h678, 12'h567, 12'h779, 12'h89a, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h89b, 12'h78a, 12'h789, 12'h679, 12'h678, 12'h679, 12'h679, 12'h678, 12'h568, 12'h467, 12'h467, 12'h568, 12'h568, 12'h578, 12'h679, 12'h89a, 12'h9ab, 12'habc, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbbe, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'habc, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h789, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'h99a, 12'h889, 12'h99a, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h778, 12'h999, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbbb, 12'h99a, 12'h899, 12'h788, 12'h678, 12'h678, 12'h568, 12'h678, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h778, 12'h789, 12'h789, 12'h789, 12'h789, 12'h689, 12'h679, 12'h678, 12'h678, 12'h679, 12'h679, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h579, 12'h679, 12'h679, 12'h578, 12'h357, 12'h357, 12'h467, 12'h568, 12'h578, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h678, 12'h568, 12'h457, 12'h457, 12'h456, 12'h446, 12'h446, 12'h345, 12'h335, 12'h345, 
12'h445, 12'h446, 12'h456, 12'h556, 12'h456, 12'h456, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h456, 12'h557, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h668, 12'h678, 12'h678, 12'h667, 12'h667, 12'h667, 12'h677, 12'h778, 12'h888, 12'haaa, 12'hbbc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccb, 12'h998, 12'h766, 12'h666, 12'h666, 12'h766, 12'h777, 12'h877, 12'h877, 12'h777, 12'h777, 12'h777, 12'h888, 12'h887, 12'h888, 12'h888, 12'h889, 12'h899, 12'h9ab, 12'habc, 12'hbce, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcde, 12'hcdf, 
12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ab, 12'h8ab, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ab, 12'h8ac, 12'h8bc, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h8ac, 12'h79b, 12'h789, 12'h678, 12'h667, 12'h667, 12'h566, 12'h566, 12'h565, 12'h666, 12'h566, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hbbc, 12'h788, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h789, 12'h89b, 12'h9bc, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bc, 12'h9ac, 12'h89b, 12'h679, 12'h568, 12'h568, 12'h678, 12'h678, 12'h578, 12'h567, 12'h467, 12'h457, 12'h357, 12'h457, 12'h467, 12'h468, 12'h568, 12'h568, 12'h679, 12'h78a, 12'h89b, 12'habd, 12'habd, 12'hbcd, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'haac, 12'habc, 12'habc, 12'haac, 12'habd, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h89b, 12'h789, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h677, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbc, 12'h889, 12'h889, 12'h889, 12'h889, 12'h89a, 12'h99b, 12'h9ab, 12'h9ac, 12'haac, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'hace, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h779, 12'h789, 12'h789, 12'h778, 12'h777, 12'h667, 12'h667, 12'h666, 12'h666, 12'h566, 12'h666, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h666, 12'h778, 12'h999, 12'hbbb, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h889, 12'h788, 12'h778, 12'h678, 12'h678, 12'h568, 12'h567, 12'h567, 12'h567, 12'h557, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h556, 12'h566, 12'h667, 12'h667, 12'h678, 12'h678, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h578, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h579, 12'h579, 12'h579, 12'h569, 12'h579, 12'h679, 12'h578, 12'h467, 12'h357, 12'h457, 12'h467, 12'h457, 12'h568, 12'h578, 12'h679, 12'h779, 12'h779, 12'h679, 12'h678, 12'h668, 12'h567, 12'h457, 12'h456, 12'h456, 12'h456, 12'h446, 12'h445, 12'h445, 
12'h446, 12'h456, 12'h556, 12'h557, 12'h557, 12'h557, 12'h456, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h456, 12'h557, 12'h557, 12'h557, 12'h567, 12'h567, 12'h667, 12'h678, 12'h678, 12'h678, 12'h678, 12'h667, 12'h667, 12'h677, 12'h777, 12'h788, 12'h99a, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h998, 12'h776, 12'h665, 12'h666, 12'h776, 12'h777, 12'h887, 12'h877, 12'h777, 12'h777, 12'h777, 12'h877, 12'h888, 12'h888, 12'h888, 12'h899, 12'h99a, 12'h9ab, 12'habc, 12'hbce, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 
12'hcde, 12'hcce, 12'hbce, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'h9ac, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h89b, 12'h89b, 12'h8ab, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h79a, 12'h79a, 12'h79a, 12'h79a, 12'h89a, 12'h79a, 12'h79a, 12'h89a, 12'h8ac, 12'h8bc, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bc, 12'h8ac, 12'h8ab, 12'h79a, 12'h678, 12'h677, 12'h667, 12'h566, 12'h666, 12'h666, 12'h566, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h99a, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h79a, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h89b, 12'h78a, 12'h468, 12'h568, 12'h568, 12'h567, 12'h567, 12'h467, 12'h467, 12'h457, 12'h457, 12'h457, 12'h467, 12'h568, 12'h568, 12'h568, 12'h679, 12'h679, 12'h78a, 12'h88a, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbd, 12'hbbd, 12'habd, 12'haac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h9ab, 12'h9ac, 12'h9ac, 12'habc, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h89a, 12'h789, 12'h577, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'h99a, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h779, 12'h889, 12'h89a, 12'h99b, 12'h9ac, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h889, 12'h789, 12'h778, 12'h678, 12'h667, 12'h667, 12'h566, 12'h566, 12'h566, 12'h666, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h565, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h555, 12'h655, 12'h666, 12'h666, 12'h667, 12'h788, 12'h999, 12'hbbb, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h99a, 12'h899, 12'h889, 12'h788, 12'h789, 12'h779, 12'h678, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h556, 12'h557, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h567, 12'h667, 12'h667, 12'h677, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h467, 12'h467, 12'h568, 12'h568, 12'h568, 12'h678, 12'h578, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h456, 12'h346, 12'h356, 12'h456, 12'h457, 12'h467, 12'h568, 12'h679, 12'h679, 12'h779, 12'h679, 12'h678, 12'h568, 12'h567, 12'h456, 12'h346, 12'h446, 12'h456, 12'h456, 12'h446, 12'h556, 
12'h456, 12'h556, 12'h557, 12'h567, 12'h667, 12'h567, 12'h557, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h678, 12'h678, 12'h678, 12'h667, 12'h667, 12'h667, 12'h677, 12'h778, 12'h999, 12'hbbb, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdcc, 12'haa9, 12'h777, 12'h666, 12'h666, 12'h666, 12'h777, 12'h887, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h99a, 12'h9aa, 12'h9ab, 12'habc, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcde, 12'hcce, 
12'hbcd, 12'hbcd, 12'hbcd, 12'hbbc, 12'habc, 12'hbbc, 12'habc, 12'habc, 12'h9ab, 12'h9ab, 12'h9ab, 12'haac, 12'h9ab, 12'h89b, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h89a, 12'h889, 12'h78a, 12'h789, 12'h778, 12'h678, 12'h678, 12'h677, 12'h677, 12'h678, 12'h788, 12'h789, 12'h789, 12'h788, 12'h788, 12'h789, 12'h79a, 12'h8ab, 12'h8bc, 12'h9bd, 12'h9bc, 12'h9bd, 12'h9bd, 12'h8bc, 12'h8ac, 12'h89b, 12'h789, 12'h677, 12'h666, 12'h555, 12'h566, 12'h666, 12'h566, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h99a, 12'h567, 12'h567, 12'h677, 12'h567, 12'h567, 12'h567, 12'h679, 12'h89b, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h78a, 12'h579, 12'h467, 12'h468, 12'h568, 12'h568, 12'h467, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h679, 12'h679, 12'h679, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbd, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h89b, 12'h89a, 12'h78a, 12'h789, 12'h789, 12'h679, 12'h679, 12'h679, 12'h789, 12'h789, 12'h679, 12'h689, 
12'h78a, 12'h89a, 12'h89b, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h89b, 12'h789, 12'h678, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h667, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h9aa, 12'h888, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h789, 12'h89b, 12'h99b, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h78a, 12'h88a, 12'h789, 12'h778, 12'h778, 12'h678, 12'h667, 12'h667, 12'h566, 12'h566, 12'h556, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h655, 12'h665, 12'h666, 12'h667, 12'h778, 12'h899, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'habb, 12'h999, 12'h889, 12'h888, 12'h889, 12'h789, 12'h788, 12'h678, 12'h567, 12'h567, 12'h678, 12'h568, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h567, 12'h667, 12'h667, 12'h667, 12'h567, 12'h567, 12'h667, 12'h567, 12'h567, 12'h467, 12'h467, 12'h557, 12'h567, 12'h568, 12'h578, 12'h578, 12'h568, 12'h568, 12'h567, 12'h567, 12'h567, 12'h467, 12'h456, 12'h346, 12'h356, 12'h356, 12'h356, 12'h457, 12'h457, 12'h568, 12'h668, 12'h679, 12'h679, 12'h668, 12'h568, 12'h567, 12'h456, 12'h346, 12'h346, 12'h446, 12'h446, 12'h446, 12'h456, 
12'h456, 12'h556, 12'h567, 12'h667, 12'h667, 12'h667, 12'h557, 12'h456, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h557, 12'h567, 12'h667, 12'h678, 12'h667, 12'h567, 12'h567, 12'h667, 12'h677, 12'h778, 12'h899, 12'haaa, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbba, 12'h888, 12'h776, 12'h666, 12'h666, 12'h777, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h887, 12'h888, 12'h899, 12'h99a, 12'h9aa, 12'h9ab, 12'habd, 12'hbce, 12'hbde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hccd, 
12'habc, 12'habc, 12'habb, 12'haab, 12'haab, 12'haab, 12'h99a, 12'h899, 12'h889, 12'h888, 12'h889, 12'h99a, 12'h9aa, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h678, 12'h667, 12'h667, 12'h566, 12'h556, 12'h556, 12'h566, 12'h566, 12'h677, 12'h678, 12'h678, 12'h678, 12'h678, 12'h789, 12'h79a, 12'h89b, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ac, 12'h79a, 12'h678, 12'h666, 12'h555, 12'h566, 12'h566, 12'h566, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haab, 12'h567, 12'h677, 12'h667, 12'h567, 12'h567, 12'h567, 12'h78a, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h89b, 12'h568, 12'h568, 12'h579, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h789, 12'h789, 12'h789, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h78b, 12'h89b, 12'h89b, 12'h9ac, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbd, 12'habd, 12'h9ac, 12'h89b, 12'h89b, 12'h78a, 12'h679, 12'h679, 12'h668, 12'h568, 12'h568, 12'h568, 12'h568, 12'h567, 12'h567, 12'h568, 12'h568, 12'h578, 
12'h679, 12'h789, 12'h789, 12'h89a, 12'h9ac, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h89b, 12'h789, 12'h678, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h889, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hccd, 12'haab, 12'h999, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h789, 12'h89a, 12'h99b, 12'h9ac, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 
12'habe, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'habe, 12'hace, 12'hace, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h789, 12'h789, 12'h778, 12'h778, 12'h667, 12'h667, 12'h666, 12'h566, 12'h555, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h565, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h777, 12'h899, 12'hbbb, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h889, 12'h888, 12'h788, 12'h788, 12'h788, 12'h678, 12'h668, 12'h678, 12'h678, 12'h568, 12'h567, 12'h568, 12'h667, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h556, 12'h556, 12'h556, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h667, 12'h567, 12'h567, 12'h567, 12'h457, 12'h457, 12'h567, 12'h567, 12'h568, 12'h568, 12'h568, 12'h568, 12'h567, 12'h467, 12'h456, 12'h456, 12'h456, 12'h346, 12'h356, 12'h355, 12'h356, 12'h457, 12'h457, 12'h457, 12'h568, 12'h668, 12'h668, 12'h568, 12'h567, 12'h467, 12'h456, 12'h346, 12'h346, 12'h446, 12'h446, 12'h446, 12'h446, 
12'h446, 12'h456, 12'h557, 12'h667, 12'h667, 12'h667, 12'h567, 12'h557, 12'h456, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h456, 12'h556, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h566, 12'h566, 12'h566, 12'h667, 12'h778, 12'h888, 12'haaa, 12'hbbb, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccb, 12'h999, 12'h777, 12'h666, 12'h666, 12'h777, 12'h887, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h877, 12'h888, 12'h899, 12'h99a, 12'h9aa, 12'h9ab, 12'hbcd, 12'hbce, 12'hbde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbcd, 12'habc, 
12'h9aa, 12'h9aa, 12'h999, 12'h999, 12'h899, 12'h888, 12'h788, 12'h778, 12'h778, 12'h889, 12'h888, 12'h788, 12'h899, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h8ab, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h788, 12'h678, 12'h677, 12'h677, 12'h667, 12'h566, 12'h566, 12'h666, 12'h567, 12'h667, 12'h667, 12'h678, 12'h778, 12'h788, 12'h789, 12'h789, 12'h89a, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h89b, 12'h789, 12'h677, 12'h566, 12'h556, 12'h566, 12'h666, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h678, 12'h678, 12'h567, 12'h567, 12'h567, 12'h578, 12'h89b, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h79b, 12'h679, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'h9ac, 12'h89b, 12'h78a, 12'h78a, 12'h679, 12'h679, 12'h669, 12'h568, 12'h568, 12'h568, 12'h567, 12'h467, 12'h467, 12'h457, 12'h457, 12'h467, 12'h467, 
12'h568, 12'h678, 12'h679, 12'h789, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h9ab, 12'h789, 12'h678, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h899, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbbb, 12'h99a, 12'h889, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h789, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'hace, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h78a, 12'h789, 12'h789, 12'h778, 12'h678, 12'h667, 12'h667, 12'h566, 12'h556, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h565, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h566, 12'h666, 12'h778, 12'h999, 12'hbbb, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h9aa, 12'h889, 12'h889, 12'h888, 12'h788, 12'h788, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h568, 12'h567, 12'h667, 12'h668, 12'h667, 12'h556, 12'h456, 12'h456, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h556, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h567, 12'h556, 12'h456, 12'h457, 12'h457, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h457, 12'h456, 12'h456, 12'h456, 12'h345, 12'h455, 12'h355, 12'h355, 12'h356, 12'h456, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h568, 12'h457, 12'h557, 12'h457, 12'h456, 12'h446, 12'h446, 12'h345, 12'h346, 12'h346, 
12'h346, 12'h446, 12'h456, 12'h557, 12'h567, 12'h567, 12'h557, 12'h556, 12'h556, 12'h456, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h446, 12'h456, 12'h567, 12'h557, 12'h557, 12'h557, 12'h456, 12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h667, 12'h778, 12'h999, 12'habb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hccc, 12'h999, 12'h777, 12'h665, 12'h776, 12'h777, 12'h887, 12'h888, 12'h777, 12'h777, 12'h776, 12'h666, 12'h777, 12'h888, 12'h899, 12'h99a, 12'h9ab, 12'h9bc, 12'hbcd, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hcde, 12'hcce, 12'hbcd, 12'habc, 12'h99a, 
12'h999, 12'h899, 12'h888, 12'h888, 12'h788, 12'h778, 12'h778, 12'h777, 12'h777, 12'h788, 12'h889, 12'h889, 12'h889, 12'h899, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h88a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h8ab, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h678, 12'h678, 12'h677, 12'h677, 12'h677, 12'h678, 12'h678, 12'h678, 12'h678, 12'h788, 12'h678, 12'h788, 12'h789, 12'h89b, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bc, 12'h8ac, 12'h79a, 12'h678, 12'h555, 12'h555, 12'h566, 12'h666, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbbc, 12'h678, 12'h677, 12'h567, 12'h567, 12'h567, 12'h678, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'hacd, 12'habd, 12'h9ac, 12'h89c, 12'h79b, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h88b, 12'h78a, 12'h67a, 12'h77a, 12'h679, 12'h679, 12'h679, 12'h678, 12'h678, 12'h568, 12'h568, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 
12'h467, 12'h567, 12'h568, 12'h678, 12'h78a, 12'h9ab, 12'haac, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h89a, 12'h679, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h9aa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'habb, 12'h99a, 12'h89a, 12'h889, 12'h889, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h677, 12'h678, 12'h778, 12'h88a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 
12'hccf, 12'hccf, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'habe, 12'habe, 12'hace, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h79b, 12'h78a, 12'h78a, 12'h78a, 12'h89a, 12'h78a, 12'h78a, 12'h789, 12'h779, 12'h678, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h667, 12'h666, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'h788, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'habb, 12'h999, 12'h888, 12'h788, 12'h778, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h568, 12'h567, 12'h667, 12'h567, 12'h567, 12'h456, 12'h445, 12'h455, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h446, 12'h446, 12'h557, 12'h667, 12'h668, 12'h668, 12'h668, 12'h677, 12'h677, 12'h677, 12'h667, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h467, 12'h567, 12'h567, 12'h567, 12'h467, 12'h457, 12'h456, 12'h456, 12'h456, 12'h345, 12'h455, 12'h455, 12'h346, 12'h356, 12'h456, 12'h457, 12'h557, 12'h568, 12'h568, 12'h568, 12'h567, 12'h457, 12'h557, 12'h557, 12'h557, 12'h456, 12'h446, 12'h346, 12'h346, 12'h346, 
12'h446, 12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h456, 12'h456, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h556, 12'h456, 12'h456, 12'h345, 12'h445, 12'h455, 12'h455, 12'h456, 12'h556, 12'h556, 12'h666, 12'h777, 12'h889, 12'haaa, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haa9, 12'h777, 12'h666, 12'h776, 12'h777, 12'h877, 12'h887, 12'h777, 12'h777, 12'h666, 12'h666, 12'h776, 12'h887, 12'h888, 12'h89a, 12'h9ab, 12'habd, 12'hbce, 12'hbde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbcd, 12'hbcd, 12'habb, 12'h99a, 12'h899, 
12'h889, 12'h888, 12'h888, 12'h778, 12'h778, 12'h788, 12'h788, 12'h788, 12'h888, 12'h889, 12'h899, 12'h99a, 12'h89a, 12'h89a, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h8ab, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h789, 12'h79a, 12'h89a, 12'h79a, 12'h89a, 12'h89a, 12'h79a, 12'h789, 12'h789, 12'h678, 12'h788, 12'h789, 12'h8ab, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h89b, 12'h688, 12'h566, 12'h555, 12'h555, 12'h566, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h678, 12'h567, 12'h567, 12'h567, 12'h567, 12'h679, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'hacd, 12'habd, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h679, 12'h578, 12'h568, 12'h457, 12'h457, 12'h457, 12'h467, 
12'h467, 12'h467, 12'h467, 12'h567, 12'h568, 12'h789, 12'h9ab, 12'haac, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h89a, 12'h789, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'habb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccd, 12'haab, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h88a, 12'h889, 12'h889, 12'h889, 12'h879, 12'h778, 12'h778, 12'h778, 12'h778, 12'h678, 12'h778, 12'h789, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79a, 12'h79a, 12'h89a, 12'h88a, 12'h88a, 12'h789, 12'h789, 12'h778, 12'h678, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h666, 12'h565, 12'h565, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h788, 12'h677, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h456, 12'h345, 12'h445, 12'h445, 12'h445, 12'h345, 12'h335, 12'h335, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h557, 12'h667, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h677, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h456, 12'h446, 12'h445, 12'h455, 12'h456, 12'h356, 12'h456, 12'h457, 12'h567, 12'h568, 12'h568, 12'h568, 12'h457, 12'h457, 12'h457, 12'h557, 12'h567, 12'h567, 12'h456, 12'h446, 12'h346, 12'h346, 
12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h456, 12'h567, 12'h567, 12'h567, 12'h667, 12'h567, 12'h556, 12'h456, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h556, 12'h556, 12'h667, 12'h778, 12'h999, 12'haab, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h877, 12'h666, 12'h766, 12'h777, 12'h887, 12'h888, 12'h777, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h888, 12'h89a, 12'h9ab, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbcd, 12'hbbc, 12'haab, 12'h9aa, 12'h999, 12'h889, 
12'h889, 12'h889, 12'h889, 12'h888, 12'h889, 12'h899, 12'h99a, 12'h99a, 12'h999, 12'h99a, 12'h9aa, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9aa, 12'h9ab, 12'h99a, 12'h89a, 12'h99b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ab, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h9ac, 12'h8ab, 12'h89b, 12'h89a, 12'h799, 12'h789, 12'h79a, 12'h8ab, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h789, 12'h566, 12'h555, 12'h555, 12'h566, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hddd, 12'h789, 12'h678, 12'h678, 12'h567, 12'h567, 12'h78a, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hacd, 12'habd, 12'h9ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbbe, 12'hbbe, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h78a, 12'h789, 12'h679, 12'h568, 12'h568, 
12'h568, 12'h568, 12'h467, 12'h467, 12'h568, 12'h679, 12'h89a, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'haac, 12'h89b, 12'h789, 12'h678, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcd, 12'habc, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h99b, 12'h89a, 12'h88a, 12'h88a, 12'h889, 12'h789, 12'h779, 12'h778, 12'h778, 12'h779, 12'h789, 12'h88a, 12'h99b, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 
12'hccf, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h89b, 12'h89a, 12'h89a, 12'h88a, 12'h889, 12'h789, 12'h778, 12'h778, 12'h777, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'h899, 12'haab, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h9aa, 12'h889, 12'h788, 12'h778, 12'h677, 12'h667, 12'h677, 12'h678, 12'h678, 12'h678, 12'h678, 12'h667, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h456, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h446, 12'h556, 12'h567, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h677, 12'h677, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h556, 12'h556, 12'h456, 12'h456, 12'h455, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h568, 12'h668, 12'h568, 12'h457, 12'h457, 12'h456, 12'h457, 12'h557, 12'h567, 12'h456, 12'h346, 12'h346, 12'h346, 
12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h345, 12'h445, 12'h446, 12'h445, 12'h445, 12'h446, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h666, 12'h566, 12'h556, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h566, 12'h777, 12'h889, 12'haaa, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedd, 12'hbbb, 12'h888, 12'h666, 12'h776, 12'h777, 12'h887, 12'h887, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h9aa, 12'habd, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'hbbc, 12'habb, 12'h9ab, 12'h99a, 12'h999, 12'h899, 
12'h99a, 12'h9aa, 12'haaa, 12'haab, 12'habb, 12'habb, 12'haab, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h89b, 12'h8ab, 12'h89b, 12'h8ab, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h89b, 12'h89b, 12'h8ab, 12'h9bc, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h79a, 12'h666, 12'h455, 12'h555, 12'h556, 12'h666, 12'h566, 12'h555, 12'h555, 12'h666, 12'h999, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h889, 12'h678, 12'h668, 12'h567, 12'h567, 12'h89b, 12'habd, 12'habd, 12'hace, 12'hace, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h89c, 12'h99c, 12'h9ac, 12'h99c, 12'h99c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h789, 
12'h779, 12'h679, 12'h568, 12'h568, 12'h457, 12'h568, 12'h78a, 12'h89b, 12'h9ac, 12'habc, 12'habc, 12'habc, 12'h9ab, 12'h89a, 12'h678, 12'h567, 12'h456, 12'h456, 12'h466, 12'h567, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hddd, 12'hccd, 12'hbcc, 12'haac, 12'h9ab, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h88a, 12'h78a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h78a, 12'h89b, 12'h9ac, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 
12'hbce, 12'hbce, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h778, 12'h777, 12'h677, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h777, 12'h999, 12'habb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h888, 12'h778, 12'h777, 12'h667, 12'h567, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h456, 12'h456, 12'h445, 12'h445, 12'h345, 12'h345, 12'h335, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h556, 12'h556, 12'h557, 12'h557, 12'h667, 12'h667, 12'h677, 12'h778, 12'h667, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h557, 12'h667, 12'h667, 12'h567, 12'h557, 12'h556, 12'h556, 12'h456, 12'h456, 12'h446, 12'h456, 12'h456, 12'h456, 12'h467, 12'h567, 12'h568, 12'h668, 12'h568, 12'h567, 12'h457, 12'h457, 12'h457, 12'h457, 12'h557, 12'h456, 12'h446, 12'h446, 12'h457, 
12'h457, 12'h457, 12'h557, 12'h557, 12'h457, 12'h457, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h556, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h556, 12'h667, 12'h778, 12'h999, 12'haab, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'hccb, 12'h999, 12'h777, 12'h776, 12'h777, 12'h887, 12'h887, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h778, 12'h899, 12'habc, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbcd, 12'habc, 12'haab, 12'h99a, 12'h99a, 12'h9aa, 12'haab, 
12'habb, 12'hbbc, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'habc, 12'habc, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9ac, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bc, 12'h89b, 12'h677, 12'h455, 12'h455, 12'h555, 12'h666, 12'h666, 12'h555, 12'h555, 12'h666, 12'h9aa, 
12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h778, 12'h678, 12'h678, 12'h567, 12'h678, 12'h9ab, 12'habd, 12'habd, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 
12'h88a, 12'h78a, 12'h679, 12'h679, 12'h568, 12'h468, 12'h679, 12'h89b, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h89b, 12'h678, 12'h567, 12'h567, 12'h456, 12'h456, 12'h677, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccd, 12'hbcc, 12'hbbc, 12'habb, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haac, 12'h9ac, 12'h89b, 12'h88b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h789, 12'h88a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'hbbd, 12'hbce, 12'hcce, 12'hcdf, 12'hddf, 12'hddf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h778, 12'h777, 12'h677, 12'h666, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h787, 12'h999, 12'hbbb, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hccc, 12'habb, 12'h999, 12'h888, 12'h778, 12'h677, 12'h567, 12'h556, 12'h566, 12'h667, 12'h667, 12'h678, 12'h677, 12'h567, 12'h567, 12'h556, 12'h556, 12'h556, 12'h556, 12'h445, 12'h445, 12'h345, 12'h335, 12'h345, 12'h335, 12'h335, 12'h345, 12'h345, 12'h445, 12'h445, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h667, 12'h667, 12'h778, 12'h778, 12'h667, 12'h667, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h667, 12'h667, 12'h668, 12'h667, 12'h667, 12'h567, 12'h456, 12'h446, 12'h446, 12'h446, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h668, 12'h678, 12'h678, 12'h668, 12'h568, 12'h568, 12'h558, 12'h557, 12'h457, 12'h457, 12'h447, 12'h557, 12'h558, 
12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h457, 12'h447, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h567, 12'h567, 12'h567, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h344, 12'h345, 12'h445, 12'h455, 12'h556, 12'h677, 12'h889, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'ha99, 12'h777, 12'h776, 12'h777, 12'h887, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h676, 12'h888, 12'h9aa, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbbc, 12'h9ab, 12'h99a, 12'h9aa, 12'haab, 12'habb, 12'hbcd, 
12'hccd, 12'hccd, 12'hbce, 12'hbce, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ab, 12'h678, 12'h555, 12'h455, 12'h566, 12'h666, 12'h666, 12'h555, 12'h555, 12'h676, 12'haaa, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h678, 12'h678, 12'h568, 12'h568, 12'h679, 12'h9ac, 12'habd, 12'habd, 12'hbce, 12'hace, 12'hace, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 
12'h89b, 12'h89b, 12'h78a, 12'h679, 12'h679, 12'h579, 12'h579, 12'h79a, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'haac, 12'h9ab, 12'h789, 12'h567, 12'h567, 12'h567, 12'h466, 12'h788, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccc, 12'hbcc, 12'hbcc, 12'habc, 12'haab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'haad, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h89b, 12'h99c, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'habd, 12'haad, 12'haac, 12'habc, 
12'habc, 12'habd, 12'habc, 12'hbbd, 12'hbce, 12'hcce, 12'hcde, 12'hcde, 12'hcce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h778, 12'h778, 12'h677, 12'h666, 12'h666, 12'h666, 12'h565, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h899, 12'h788, 12'h777, 12'h667, 12'h556, 12'h556, 12'h566, 12'h667, 12'h667, 12'h678, 12'h678, 12'h667, 12'h566, 12'h556, 12'h556, 12'h556, 12'h456, 12'h445, 12'h345, 12'h345, 12'h335, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h445, 12'h445, 12'h445, 12'h455, 12'h556, 12'h556, 12'h556, 12'h667, 12'h778, 12'h778, 12'h778, 12'h667, 12'h567, 12'h556, 12'h456, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h567, 12'h667, 12'h678, 12'h778, 12'h778, 12'h677, 12'h667, 12'h556, 12'h456, 12'h446, 12'h446, 12'h456, 12'h456, 12'h567, 12'h567, 12'h568, 12'h678, 12'h679, 12'h679, 12'h77a, 12'h77a, 12'h679, 12'h669, 12'h558, 12'h458, 12'h458, 12'h558, 12'h568, 12'h569, 
12'h569, 12'h669, 12'h669, 12'h679, 12'h568, 12'h458, 12'h357, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h556, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h456, 12'h556, 12'h556, 12'h456, 12'h445, 12'h445, 12'h345, 12'h344, 12'h334, 12'h344, 12'h334, 12'h345, 12'h445, 12'h455, 12'h667, 12'h778, 12'h99a, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbba, 12'h998, 12'h777, 12'h776, 12'h777, 12'h887, 12'h777, 12'h666, 12'h666, 12'h555, 12'h666, 12'h777, 12'h999, 12'habc, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'haab, 12'h9ab, 12'haab, 12'habc, 12'hbcd, 12'hcde, 12'hcde, 
12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ab, 12'h678, 12'h555, 12'h455, 12'h556, 12'h666, 12'h566, 12'h555, 12'h555, 12'h677, 12'haaa, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'h99a, 12'h678, 12'h678, 12'h678, 12'h678, 12'h789, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h9ac, 12'habc, 12'habc, 12'habd, 12'habc, 12'h9ab, 12'h789, 12'h567, 12'h567, 12'h567, 12'h567, 12'h99a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'hddd, 12'hbcc, 12'habb, 12'hbcc, 12'hbbc, 12'habc, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ab, 12'h99b, 12'h89b, 12'h99b, 12'h9ab, 12'haac, 12'hbbd, 12'hbbd, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h789, 12'h778, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h565, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h778, 12'h677, 12'h666, 12'h556, 12'h556, 12'h556, 12'h667, 12'h667, 12'h677, 12'h677, 12'h667, 12'h566, 12'h556, 12'h456, 12'h556, 12'h456, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h345, 12'h445, 12'h445, 12'h445, 12'h456, 12'h556, 12'h566, 12'h778, 12'h888, 12'h788, 12'h678, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h556, 12'h567, 12'h677, 12'h678, 12'h778, 12'h778, 12'h677, 12'h667, 12'h556, 12'h456, 12'h446, 12'h446, 12'h456, 12'h557, 12'h567, 12'h568, 12'h668, 12'h679, 12'h78a, 12'h78b, 12'h88b, 12'h88b, 12'h78b, 12'h67a, 12'h56a, 12'h569, 12'h569, 12'h66a, 12'h67a, 12'h67a, 
12'h57a, 12'h67a, 12'h67a, 12'h67a, 12'h679, 12'h568, 12'h357, 12'h347, 12'h447, 12'h446, 12'h446, 12'h446, 12'h556, 12'h556, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h556, 12'h456, 12'h445, 12'h445, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h445, 12'h556, 12'h777, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haa9, 12'h888, 12'h777, 12'h777, 12'h777, 12'h887, 12'h777, 12'h666, 12'h565, 12'h565, 12'h666, 12'h888, 12'h9aa, 12'hbbc, 12'hcde, 12'hcdf, 12'hcde, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hbcd, 12'habc, 12'habc, 12'hbbc, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 
12'hcde, 12'hcce, 12'hbce, 12'hbce, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ab, 12'h678, 12'h555, 12'h455, 12'h555, 12'h666, 12'h566, 12'h555, 12'h555, 12'h777, 12'haaa, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h889, 12'h89a, 12'h78a, 12'h578, 12'h678, 12'h89a, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h9ac, 12'haac, 12'habc, 12'habd, 12'habc, 12'h9ac, 12'h78a, 12'h568, 12'h567, 12'h567, 12'h567, 12'habb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hccd, 12'hbbc, 12'habb, 12'habb, 12'hbbc, 12'hbbc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'habd, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 
12'h88a, 12'h889, 12'h789, 12'h789, 12'h789, 12'h789, 12'h88a, 12'h99b, 12'haac, 12'habc, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h778, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h777, 12'h899, 12'haaa, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'haaa, 12'h888, 12'h778, 12'h667, 12'h556, 12'h455, 12'h556, 12'h556, 12'h667, 12'h667, 12'h677, 12'h667, 12'h567, 12'h566, 12'h556, 12'h456, 12'h556, 12'h556, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h334, 12'h334, 12'h345, 12'h445, 12'h445, 12'h445, 12'h446, 12'h556, 12'h567, 12'h778, 12'h789, 12'h788, 12'h667, 12'h567, 12'h567, 12'h567, 12'h457, 12'h457, 12'h457, 12'h457, 12'h557, 12'h567, 12'h567, 12'h567, 12'h667, 12'h677, 12'h677, 12'h677, 12'h667, 12'h556, 12'h556, 12'h556, 12'h456, 12'h556, 12'h557, 12'h568, 12'h568, 12'h679, 12'h68a, 12'h78b, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h78b, 12'h67b, 12'h67a, 12'h68b, 12'h78b, 12'h78b, 12'h78b, 
12'h68b, 12'h67a, 12'h67a, 12'h67a, 12'h67a, 12'h569, 12'h458, 12'h347, 12'h457, 12'h457, 12'h446, 12'h456, 12'h556, 12'h556, 12'h667, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h345, 12'h445, 12'h556, 12'h667, 12'h889, 12'haab, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccb, 12'h999, 12'h887, 12'h777, 12'h777, 12'h777, 12'h887, 12'h777, 12'h666, 12'h666, 12'h665, 12'h666, 12'h888, 12'h9ab, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hbcd, 12'hbbd, 12'hbcd, 12'hccd, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hcde, 12'hbce, 12'hbce, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h788, 12'h565, 12'h555, 12'h556, 12'h566, 12'h666, 12'h555, 12'h555, 12'h777, 12'haaa, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hbbc, 12'habc, 12'habd, 12'h89b, 12'h679, 12'h679, 12'h89b, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habc, 12'h88a, 12'h568, 12'h567, 12'h567, 12'h567, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbcc, 12'hbbb, 12'habb, 12'habb, 12'haab, 12'h9aa, 12'hbbb, 12'hbbc, 12'hbbc, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 
12'h789, 12'h778, 12'h778, 12'h778, 12'h678, 12'h678, 12'h778, 12'h779, 12'h789, 12'h89a, 12'h9ab, 12'haac, 12'haac, 12'habc, 12'haac, 12'haad, 12'habd, 12'haad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h78a, 12'h789, 12'h789, 12'h778, 12'h778, 12'h677, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'h667, 12'h556, 12'h455, 12'h556, 12'h556, 12'h667, 12'h667, 12'h777, 12'h667, 12'h567, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h445, 12'h344, 12'h334, 12'h334, 12'h334, 12'h344, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h567, 12'h678, 12'h779, 12'h778, 12'h678, 12'h567, 12'h568, 12'h568, 12'h568, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h566, 12'h667, 12'h667, 12'h667, 12'h556, 12'h556, 12'h456, 12'h556, 12'h567, 12'h568, 12'h568, 12'h579, 12'h67a, 12'h78b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 
12'h68b, 12'h68b, 12'h68b, 12'h68b, 12'h67a, 12'h57a, 12'h569, 12'h458, 12'h457, 12'h557, 12'h556, 12'h456, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h556, 12'h556, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h345, 12'h445, 12'h456, 12'h667, 12'h888, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'ha99, 12'h887, 12'h777, 12'h777, 12'h777, 12'h887, 12'h777, 12'h666, 12'h665, 12'h666, 12'h666, 12'h888, 12'h9ab, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hddf, 12'hddf, 12'hcde, 12'hcde, 
12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'h9cd, 12'h9cd, 12'h9bd, 12'h9bc, 12'h789, 12'h566, 12'h555, 12'h556, 12'h666, 12'h566, 12'h555, 12'h555, 12'h677, 12'hbbb, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbcd, 12'h9ad, 12'h89c, 12'h89b, 12'h679, 12'h679, 12'h9ac, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h78a, 12'h67a, 12'h679, 12'h679, 12'h679, 12'h578, 12'h578, 12'h689, 12'h78a, 12'h89a, 12'h89b, 12'h78b, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habc, 12'h88a, 12'h568, 12'h567, 12'h567, 12'h678, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdde, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'haab, 12'haaa, 12'h99a, 12'h99a, 12'habb, 12'hbbc, 12'hbbc, 12'haab, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'h9ac, 12'habc, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 
12'h789, 12'h778, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h789, 12'h89a, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'haac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h78a, 12'h789, 12'h789, 12'h778, 12'h778, 12'h777, 12'h666, 12'h666, 12'h556, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h554, 12'h555, 12'h554, 12'h554, 12'h554, 12'h554, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'h666, 12'h556, 12'h455, 12'h455, 12'h556, 12'h666, 12'h667, 12'h777, 12'h667, 12'h567, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h445, 12'h344, 12'h334, 12'h344, 12'h334, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h567, 12'h668, 12'h679, 12'h679, 12'h679, 12'h678, 12'h679, 12'h779, 12'h789, 12'h779, 12'h678, 12'h678, 12'h567, 12'h667, 12'h567, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h567, 12'h556, 12'h556, 12'h556, 12'h556, 12'h567, 12'h678, 12'h679, 12'h579, 12'h67a, 12'h89b, 12'h9ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 
12'h79c, 12'h69c, 12'h68b, 12'h68b, 12'h68b, 12'h67a, 12'h569, 12'h468, 12'h568, 12'h568, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h456, 12'h556, 12'h556, 12'h445, 12'h445, 12'h345, 12'h445, 12'h445, 12'h445, 12'h345, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h455, 12'h666, 12'h888, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h998, 12'h877, 12'h777, 12'h777, 12'h887, 12'h777, 12'h666, 12'h555, 12'h665, 12'h666, 12'h888, 12'haab, 12'hbcd, 12'hcde, 12'hcdf, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 
12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'h9cd, 12'h9bd, 12'h9bd, 12'h799, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h555, 12'h555, 12'h777, 12'hbbc, 
12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccd, 12'h89c, 12'h78b, 12'h78b, 12'h679, 12'h68a, 12'h9ac, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'h9ac, 12'h89c, 12'h78b, 12'h57a, 12'h469, 12'h458, 12'h579, 12'h679, 12'h679, 12'h457, 12'h357, 12'h467, 12'h467, 12'h467, 12'h468, 12'h679, 12'h679, 12'h78a, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'habd, 12'habc, 12'h89a, 12'h678, 12'h567, 12'h567, 12'h789, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hccc, 12'hbbc, 12'habb, 12'haab, 12'haab, 12'h9aa, 12'h99a, 12'h778, 12'h457, 12'h346, 12'h568, 12'h679, 12'h789, 12'h88a, 12'h9ab, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 
12'h789, 12'h789, 12'h788, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h889, 12'h89a, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h889, 12'h789, 12'h889, 12'h778, 12'h778, 12'h777, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h554, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h776, 12'h888, 12'h999, 12'haab, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h666, 12'h555, 12'h445, 12'h445, 12'h445, 12'h556, 12'h667, 12'h677, 12'h667, 12'h567, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h445, 12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h446, 12'h557, 12'h667, 12'h668, 12'h679, 12'h789, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h78a, 12'h789, 12'h779, 12'h678, 12'h678, 12'h567, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h567, 12'h567, 12'h667, 12'h678, 12'h679, 12'h679, 12'h68a, 12'h89c, 12'h9ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h7ac, 12'h7ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 
12'h79d, 12'h79c, 12'h79c, 12'h78b, 12'h78b, 12'h67a, 12'h57a, 12'h569, 12'h568, 12'h668, 12'h668, 12'h668, 12'h567, 12'h567, 12'h567, 12'h557, 12'h556, 12'h556, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h445, 12'h345, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h455, 12'h666, 12'h778, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h888, 12'h887, 12'h888, 12'h887, 12'h777, 12'h666, 12'h565, 12'h666, 12'h666, 12'h788, 12'habb, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'h9cd, 12'h9bd, 12'h9bd, 12'h89a, 12'h566, 12'h556, 12'h566, 12'h566, 12'h555, 12'h555, 12'h566, 12'h789, 12'hccc, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbcd, 12'h78c, 12'h78c, 12'h78b, 12'h67a, 12'h78a, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'hbce, 12'habe, 12'habd, 12'habd, 12'h9ac, 12'h89c, 12'h79b, 12'h67a, 12'h569, 12'h569, 12'h89b, 12'haac, 12'h9ab, 12'h457, 12'h357, 12'h356, 12'h356, 12'h356, 12'h357, 12'h679, 12'h679, 12'h569, 12'h67a, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ad, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'habe, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habc, 12'habd, 12'habd, 12'habd, 12'habc, 12'h89b, 12'h678, 12'h567, 12'h678, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'hbbb, 12'hbbb, 12'hccc, 12'hcdd, 12'hddd, 12'hbbc, 12'haaa, 12'h9aa, 12'h9aa, 12'hbbb, 12'haab, 12'h889, 12'h778, 12'h778, 12'h777, 12'h667, 12'h567, 12'h678, 12'h89a, 12'habc, 12'habc, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 
12'h88a, 12'h88a, 12'h889, 12'h789, 12'h778, 12'h778, 12'h778, 12'h778, 12'h678, 12'h677, 12'h677, 12'h678, 12'h778, 12'h789, 12'h88a, 12'h89a, 12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88a, 12'h889, 12'h889, 12'h789, 12'h789, 12'h778, 12'h778, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h998, 12'h888, 12'h777, 12'h666, 12'h555, 12'h445, 12'h445, 12'h445, 12'h556, 12'h667, 12'h777, 12'h677, 12'h667, 12'h566, 12'h566, 12'h666, 12'h566, 12'h556, 12'h445, 12'h344, 12'h334, 12'h334, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h556, 12'h556, 12'h557, 12'h567, 12'h678, 12'h779, 12'h78a, 12'h78a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h78a, 12'h779, 12'h678, 12'h678, 12'h667, 12'h567, 12'h456, 12'h456, 12'h446, 12'h556, 12'h556, 12'h556, 12'h667, 12'h667, 12'h557, 12'h567, 12'h667, 12'h678, 12'h668, 12'h678, 12'h679, 12'h67a, 12'h78a, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h7ac, 12'h7ad, 12'h8ad, 12'h79d, 12'h79d, 12'h8ad, 
12'h7ad, 12'h79d, 12'h79c, 12'h79c, 12'h78b, 12'h78b, 12'h67a, 12'h679, 12'h679, 12'h679, 12'h678, 12'h668, 12'h668, 12'h668, 12'h667, 12'h567, 12'h557, 12'h556, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h244, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h345, 12'h445, 12'h556, 12'h777, 12'h899, 12'haab, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'haa9, 12'ha98, 12'h888, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h888, 12'habb, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hacd, 12'h9cd, 12'h9cd, 12'h9bd, 12'h8ab, 12'h677, 12'h556, 12'h566, 12'h566, 12'h555, 12'h566, 12'h677, 12'h89a, 12'hccd, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbd, 12'h78c, 12'h78c, 12'h78b, 12'h78a, 12'h89b, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h78b, 12'h78a, 12'h89a, 12'h9ac, 12'h9ab, 12'h568, 12'h457, 12'h246, 12'h246, 12'h246, 12'h568, 12'h89a, 12'h89a, 12'h679, 12'h458, 12'h89b, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ab, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 
12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h99b, 12'h678, 12'h567, 12'h678, 12'hbcc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'hcdd, 12'hddd, 12'hccc, 12'haab, 12'hbbb, 12'hccc, 12'hbbb, 12'h889, 12'hbbb, 12'hbbb, 12'haaa, 12'h99a, 12'h99a, 12'h99a, 12'haaa, 12'hddd, 12'hddd, 12'h999, 12'h888, 12'h666, 12'h666, 12'h555, 12'h566, 12'h89a, 12'haac, 12'haac, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 
12'h89b, 12'h89a, 12'h89a, 12'h889, 12'h789, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h788, 12'h789, 12'h789, 12'h778, 12'h779, 12'h789, 12'h88a, 12'h89a, 12'h89b, 12'h89b, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89a, 12'h89a, 12'h889, 12'h889, 12'h789, 12'h788, 12'h778, 12'h778, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h676, 12'h777, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hbbb, 12'ha99, 12'h888, 12'h888, 12'h777, 12'h566, 12'h455, 12'h445, 12'h445, 12'h445, 12'h456, 12'h667, 12'h778, 12'h777, 12'h666, 12'h556, 12'h566, 12'h667, 12'h667, 12'h556, 12'h445, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h557, 12'h557, 12'h668, 12'h678, 12'h779, 12'h789, 12'h78a, 12'h79a, 12'h89a, 12'h89a, 12'h78a, 12'h789, 12'h678, 12'h668, 12'h567, 12'h556, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h556, 12'h557, 12'h667, 12'h667, 12'h557, 12'h667, 12'h778, 12'h789, 12'h778, 12'h679, 12'h679, 12'h67a, 12'h78b, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ad, 12'h7ad, 12'h7ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 
12'h7ad, 12'h79d, 12'h89d, 12'h79c, 12'h79c, 12'h78b, 12'h67a, 12'h67a, 12'h679, 12'h679, 12'h679, 12'h678, 12'h668, 12'h678, 12'h668, 12'h667, 12'h567, 12'h557, 12'h556, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h556, 12'h667, 12'h888, 12'haaa, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'hddd, 12'hcbb, 12'hba9, 12'h998, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h888, 12'h9ab, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'hace, 12'habd, 12'habd, 
12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'h9cd, 12'h9cd, 12'h9cd, 12'h8ac, 12'h678, 12'h566, 12'h566, 12'h666, 12'h566, 12'h567, 12'h679, 12'h89b, 12'hcdd, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbd, 12'h78c, 12'h78c, 12'h89c, 12'h78b, 12'h89c, 12'habd, 12'habd, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h789, 12'h467, 12'h357, 12'h357, 12'h247, 12'h679, 12'h99b, 12'h99b, 12'h67a, 12'h469, 12'h89c, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h9ac, 12'h78b, 12'h679, 12'h679, 12'h679, 12'h568, 12'h568, 12'h568, 12'h568, 12'h679, 12'h679, 12'h78a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h9ab, 12'h679, 12'h567, 12'h688, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'heee, 12'hccd, 12'haab, 12'haaa, 12'hbbc, 12'haaa, 12'h456, 12'h778, 12'h99a, 12'h99a, 12'h999, 12'h888, 12'h777, 12'h777, 12'hbbb, 12'hccc, 12'h999, 12'h888, 12'h777, 12'h777, 12'h666, 12'h455, 12'h456, 12'h88a, 12'h9ac, 12'haac, 12'h9ac, 12'h9ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h89a, 12'h89a, 12'h889, 12'h889, 12'h889, 12'h889, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h88a, 12'h89b, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88a, 12'h889, 12'h889, 12'h889, 12'h788, 12'h778, 12'h778, 12'h778, 12'h777, 12'h666, 12'h666, 12'h666, 12'h665, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h777, 12'h888, 12'h999, 12'haab, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h888, 12'h888, 12'h777, 12'h666, 12'h455, 12'h445, 12'h445, 12'h445, 12'h455, 12'h667, 12'h778, 12'h777, 12'h666, 12'h556, 12'h566, 12'h667, 12'h667, 12'h556, 12'h445, 12'h334, 12'h334, 12'h344, 12'h344, 12'h445, 12'h445, 12'h345, 12'h345, 12'h446, 12'h456, 12'h557, 12'h557, 12'h668, 12'h668, 12'h679, 12'h679, 12'h789, 12'h78a, 12'h78a, 12'h789, 12'h779, 12'h678, 12'h668, 12'h567, 12'h556, 12'h456, 12'h445, 12'h345, 12'h446, 12'h446, 12'h446, 12'h557, 12'h667, 12'h667, 12'h667, 12'h567, 12'h668, 12'h779, 12'h789, 12'h779, 12'h679, 12'h679, 12'h67a, 12'h78b, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 
12'h79d, 12'h79d, 12'h89d, 12'h79d, 12'h79c, 12'h78b, 12'h68b, 12'h67a, 12'h67a, 12'h67a, 12'h679, 12'h679, 12'h669, 12'h678, 12'h668, 12'h568, 12'h567, 12'h567, 12'h457, 12'h456, 12'h446, 12'h446, 12'h445, 12'h345, 12'h345, 12'h345, 12'h344, 12'h334, 12'h334, 12'h234, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h445, 12'h566, 12'h777, 12'h999, 12'hbbb, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdcc, 12'hbaa, 12'h998, 12'h877, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h9aa, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'hace, 12'h9cd, 12'h9ce, 12'h9bc, 12'h688, 12'h566, 12'h666, 12'h667, 12'h567, 12'h668, 12'h78a, 12'haac, 12'hdee, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbbd, 12'h89c, 12'h78c, 12'h9ad, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89a, 12'h78a, 12'h78a, 12'h89b, 12'h9ab, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ac, 12'haad, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h569, 12'h679, 12'h78a, 12'h678, 12'h567, 12'h567, 12'h457, 12'h357, 12'h457, 12'h679, 12'h88a, 12'h679, 12'h679, 12'h679, 12'h78a, 
12'h78b, 12'h89b, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ab, 12'h679, 12'h578, 12'h9ab, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hdde, 12'hfff, 12'hdde, 12'hccc, 12'hbbb, 12'haab, 12'h888, 12'h556, 12'h556, 12'h778, 12'h99a, 12'h99a, 12'h889, 12'h788, 12'h889, 12'haab, 12'hbbb, 12'h999, 12'h778, 12'h788, 12'h888, 12'h888, 12'h788, 12'h456, 12'h457, 12'h99b, 12'haac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h99b, 12'h88a, 12'h789, 12'h779, 12'h789, 12'h889, 12'h889, 12'h789, 12'h789, 12'h88a, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89a, 12'h889, 12'h889, 12'h889, 12'h889, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h554, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h777, 12'h889, 12'haaa, 12'hbbc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hbbb, 12'h998, 12'h888, 12'h888, 12'h777, 12'h666, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h667, 12'h667, 12'h666, 12'h556, 12'h556, 12'h667, 12'h667, 12'h556, 12'h445, 12'h334, 12'h334, 12'h345, 12'h445, 12'h445, 12'h445, 12'h456, 12'h457, 12'h457, 12'h457, 12'h568, 12'h568, 12'h569, 12'h679, 12'h679, 12'h679, 12'h679, 12'h779, 12'h779, 12'h679, 12'h678, 12'h568, 12'h567, 12'h457, 12'h456, 12'h446, 12'h446, 12'h345, 12'h456, 12'h557, 12'h557, 12'h667, 12'h667, 12'h667, 12'h567, 12'h568, 12'h678, 12'h779, 12'h679, 12'h679, 12'h779, 12'h679, 12'h67a, 12'h78b, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 
12'h7ad, 12'h7ad, 12'h7ad, 12'h79d, 12'h79c, 12'h78c, 12'h68b, 12'h68b, 12'h67a, 12'h67a, 12'h67a, 12'h679, 12'h679, 12'h679, 12'h679, 12'h579, 12'h568, 12'h567, 12'h557, 12'h557, 12'h456, 12'h456, 12'h445, 12'h445, 12'h445, 12'h445, 12'h344, 12'h334, 12'h334, 12'h234, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h444, 12'h555, 12'h677, 12'h889, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddc, 12'hbaa, 12'h998, 12'h887, 12'h666, 12'h666, 12'h666, 12'h666, 12'h778, 12'h9aa, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 
12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h678, 12'h677, 12'h667, 12'h678, 12'h678, 12'h678, 12'h689, 12'h78a, 12'h79a, 12'h79b, 12'h79b, 12'h79c, 12'h7ac, 12'h8ac, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hace, 12'hace, 12'hace, 12'h9ce, 12'h9bd, 12'h789, 12'h667, 12'h666, 12'h667, 12'h678, 12'h679, 12'h89b, 12'hccd, 12'heef, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hbbd, 12'h89c, 12'h89c, 12'habd, 12'h9ad, 12'h9ad, 12'habd, 12'habe, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ad, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hccf, 12'hcdf, 12'hcdf, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'haad, 12'h89c, 12'h579, 12'h78a, 12'h89b, 12'h678, 12'h457, 12'h356, 12'h356, 12'h456, 12'h457, 12'h789, 12'h9ab, 12'h89a, 12'h679, 12'h579, 12'h569, 
12'h67a, 12'h78b, 12'h89b, 12'h89c, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ab, 12'h689, 12'h679, 12'h99b, 12'hbcd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccd, 12'heef, 12'hfff, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbb, 12'h899, 12'h678, 12'h889, 12'h9ab, 12'h9ab, 12'haab, 12'h9ab, 12'h99a, 12'haab, 12'haab, 12'h88a, 12'h668, 12'h567, 12'h667, 12'h778, 12'h899, 12'h889, 12'h668, 12'h89a, 12'habc, 12'h9ac, 12'h9ac, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'haac, 12'h9ab, 12'h89a, 12'h88a, 12'h89a, 12'h88a, 12'h889, 12'h789, 12'h789, 12'h88a, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88a, 12'h889, 12'h889, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h676, 12'h888, 12'h999, 12'haab, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hccc, 12'h998, 12'h888, 12'h888, 12'h777, 12'h666, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h667, 12'h667, 12'h556, 12'h556, 12'h556, 12'h666, 12'h667, 12'h566, 12'h445, 12'h334, 12'h334, 12'h345, 12'h345, 12'h456, 12'h557, 12'h568, 12'h568, 12'h569, 12'h569, 12'h679, 12'h679, 12'h67a, 12'h67a, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h568, 12'h568, 12'h457, 12'h457, 12'h457, 12'h447, 12'h447, 12'h447, 12'h457, 12'h557, 12'h567, 12'h667, 12'h668, 12'h668, 12'h568, 12'h568, 12'h679, 12'h789, 12'h679, 12'h679, 12'h679, 12'h679, 12'h579, 12'h67a, 12'h78b, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 
12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h79c, 12'h69c, 12'h68c, 12'h68b, 12'h68b, 12'h68b, 12'h67b, 12'h68a, 12'h68a, 12'h67a, 12'h67a, 12'h679, 12'h569, 12'h568, 12'h568, 12'h557, 12'h557, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h334, 12'h334, 12'h234, 12'h234, 12'h334, 12'h224, 12'h224, 12'h234, 12'h234, 12'h334, 12'h455, 12'h566, 12'h788, 12'h99a, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hddd, 12'hbba, 12'h998, 12'h877, 12'h666, 12'h666, 12'h665, 12'h666, 12'h788, 12'h9ab, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 
12'habd, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h89b, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'hbcd, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h679, 12'h789, 12'h789, 12'h888, 12'h777, 12'h555, 12'h566, 12'h555, 12'h556, 12'h666, 12'h778, 12'h678, 12'h667, 12'h668, 12'h68a, 12'h78a, 12'h79b, 12'h79b, 12'h7ac, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'hace, 12'hace, 12'h9ce, 12'h9ce, 12'h9bd, 12'h799, 12'h566, 12'h567, 12'h678, 12'h679, 12'h78a, 12'habc, 12'hdee, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbe, 12'h9ad, 12'h9ad, 12'habe, 12'habd, 12'h9ad, 12'habd, 12'habd, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ad, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h89b, 12'h99b, 12'h789, 12'h457, 12'h357, 12'h357, 12'h457, 12'h567, 12'h89a, 12'haab, 12'h89b, 12'h78a, 12'h679, 12'h67a, 
12'h67a, 12'h79b, 12'h89c, 12'h89c, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h689, 12'h78a, 12'h9ac, 12'haac, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hdcd, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hbcc, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'haab, 12'habc, 12'haab, 12'h99b, 12'h89a, 12'h88a, 12'h88a, 12'h789, 12'h789, 12'h778, 12'h778, 12'h889, 12'h789, 12'h89a, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 
12'habd, 12'habd, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'haac, 12'haac, 12'h9ab, 12'h99b, 12'h99a, 12'h88a, 12'h789, 12'h779, 12'h779, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88a, 12'h889, 12'h789, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h566, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h565, 12'h666, 12'h777, 12'h888, 12'h99a, 12'hbcc, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heed, 12'hccc, 12'h999, 12'h888, 12'h888, 12'h777, 12'h566, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h556, 12'h666, 12'h566, 12'h556, 12'h556, 12'h556, 12'h667, 12'h556, 12'h455, 12'h344, 12'h344, 12'h234, 12'h345, 12'h556, 12'h568, 12'h679, 12'h679, 12'h77a, 12'h68a, 12'h78a, 12'h78a, 12'h78b, 12'h78b, 12'h78b, 12'h78a, 12'h78a, 12'h77a, 12'h679, 12'h669, 12'h568, 12'h458, 12'h458, 12'h458, 12'h458, 12'h568, 12'h568, 12'h568, 12'h678, 12'h568, 12'h668, 12'h568, 12'h568, 12'h568, 12'h679, 12'h78a, 12'h89a, 12'h67a, 12'h579, 12'h579, 12'h569, 12'h569, 12'h67a, 12'h79c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h7ae, 12'h7ae, 12'h7ae, 12'h7ae, 
12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h79d, 12'h69c, 12'h69c, 12'h68c, 12'h58b, 12'h68b, 12'h68b, 12'h68b, 12'h68b, 12'h68a, 12'h68a, 12'h67a, 12'h579, 12'h569, 12'h568, 12'h568, 12'h557, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h334, 12'h234, 12'h234, 12'h234, 12'h224, 12'h224, 12'h224, 12'h234, 12'h234, 12'h334, 12'h445, 12'h556, 12'h777, 12'h899, 12'haab, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h999, 12'h877, 12'h666, 12'h666, 12'h666, 12'h666, 12'h778, 12'h9aa, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbde, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 
12'habd, 12'h9ac, 12'h9ac, 12'h89b, 12'h89a, 12'h789, 12'h789, 12'h778, 12'h677, 12'h566, 12'h566, 12'h567, 12'h667, 12'h678, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'hbbd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h78a, 12'h678, 12'h899, 12'h999, 12'h677, 12'h566, 12'h566, 12'h666, 12'h555, 12'h566, 12'h778, 12'h99a, 12'h89a, 12'h678, 12'h678, 12'h678, 12'h679, 12'h78b, 12'h79b, 12'h7ac, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9cd, 12'hace, 12'hace, 12'h9ce, 12'h9ce, 12'h9bd, 12'h79a, 12'h567, 12'h567, 12'h79a, 12'h79a, 12'h89b, 12'hccd, 12'heef, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbe, 12'haad, 12'haad, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hcce, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h89b, 12'h679, 12'h568, 12'h568, 12'h789, 12'h89a, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h78b, 
12'h89b, 12'h89c, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h78a, 12'h89b, 12'h89c, 12'h99c, 12'haad, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hccd, 12'hbcc, 12'hccd, 12'hbcd, 12'habc, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'habb, 12'habc, 12'haac, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'haab, 12'h9ab, 12'h99b, 12'h88a, 12'h88a, 12'h88a, 12'h89b, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habe, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 
12'habd, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habc, 12'habc, 12'haac, 12'h99b, 12'h99b, 12'h99a, 12'h88a, 12'h789, 12'h789, 12'h779, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89a, 12'h88a, 12'h889, 12'h789, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h776, 12'h887, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hddc, 12'haa9, 12'h888, 12'h888, 12'h777, 12'h666, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h555, 12'h455, 12'h344, 12'h344, 12'h244, 12'h345, 12'h556, 12'h678, 12'h779, 12'h68a, 12'h78a, 12'h78b, 12'h78b, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h78a, 12'h67a, 12'h67a, 12'h67a, 12'h67a, 12'h67a, 12'h67a, 12'h67a, 12'h679, 12'h779, 12'h679, 12'h669, 12'h569, 12'h569, 12'h669, 12'h78a, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h579, 12'h569, 12'h569, 12'h56a, 12'h68b, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h7ae, 12'h7ae, 12'h7ae, 
12'h7ae, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h69c, 12'h69c, 12'h68c, 12'h68b, 12'h58b, 12'h68b, 12'h68b, 12'h58b, 12'h68b, 12'h68b, 12'h67a, 12'h569, 12'h569, 12'h568, 12'h557, 12'h446, 12'h446, 12'h445, 12'h445, 12'h444, 12'h344, 12'h344, 12'h344, 12'h334, 12'h234, 12'h224, 12'h224, 12'h224, 12'h234, 12'h234, 12'h344, 12'h444, 12'h555, 12'h667, 12'h888, 12'h99a, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'hcbb, 12'h999, 12'h877, 12'h666, 12'h666, 12'h666, 12'h666, 12'h788, 12'h9aa, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbde, 12'hbce, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 
12'h89b, 12'h79b, 12'h78a, 12'h679, 12'h778, 12'h888, 12'h888, 12'h666, 12'h777, 12'h666, 12'h666, 12'h666, 12'h555, 12'h556, 12'h678, 12'h779, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcde, 12'hcce, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h789, 12'h789, 12'haaa, 12'haaa, 12'h777, 12'h555, 12'h556, 12'h455, 12'h556, 12'h566, 12'h889, 12'h9ab, 12'h89a, 12'h789, 12'h789, 12'h78a, 12'h79b, 12'h79b, 12'h8ac, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'hace, 12'hace, 12'hace, 12'h9cd, 12'h9bd, 12'h89b, 12'h567, 12'h577, 12'h89b, 12'h9bd, 12'habc, 12'hdde, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbbe, 12'h9ad, 12'haad, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'h9ad, 12'h89c, 12'h89c, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h89c, 12'h9ac, 12'habd, 12'hbce, 12'hbce, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 
12'h89c, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h78a, 12'h78b, 12'h78b, 12'h78b, 12'h99c, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hddd, 12'hccd, 12'hccd, 12'hccd, 12'hbcd, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ab, 12'haab, 12'haab, 12'h9ab, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'habc, 12'h789, 12'h779, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'habd, 12'hbbd, 12'hbbe, 12'hbbe, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 
12'habd, 12'habd, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'haac, 12'haac, 12'h9ab, 12'h99b, 12'h89a, 12'h88a, 12'h88a, 12'h789, 12'h789, 12'h88a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h89a, 12'h88a, 12'h889, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h777, 12'h888, 12'ha9a, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hddd, 12'hbba, 12'h888, 12'h888, 12'h777, 12'h667, 12'h555, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h566, 12'h666, 12'h556, 12'h556, 12'h556, 12'h455, 12'h455, 12'h455, 12'h344, 12'h344, 12'h344, 12'h345, 12'h457, 12'h678, 12'h789, 12'h68a, 12'h68a, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h77a, 12'h669, 12'h569, 12'h679, 12'h78a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h67a, 12'h569, 12'h56a, 12'h56a, 12'h78c, 12'h89d, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h7be, 
12'h7ae, 12'h7ae, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h79d, 12'h69c, 12'h69c, 12'h68c, 12'h68c, 12'h68b, 12'h68b, 12'h58b, 12'h68b, 12'h68b, 12'h67a, 12'h57a, 12'h579, 12'h569, 12'h568, 12'h457, 12'h346, 12'h345, 12'h445, 12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h234, 12'h234, 12'h234, 12'h334, 12'h234, 12'h334, 12'h345, 12'h345, 12'h445, 12'h556, 12'h778, 12'h889, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccb, 12'h999, 12'h877, 12'h766, 12'h666, 12'h666, 12'h677, 12'h778, 12'h99a, 12'hacd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'habd, 12'h9ad, 12'h9ac, 12'h89b, 
12'h78a, 12'h679, 12'h678, 12'h788, 12'haaa, 12'hbbb, 12'haaa, 12'h666, 12'h677, 12'h666, 12'h666, 12'h666, 12'h555, 12'h666, 12'h788, 12'h778, 12'h779, 12'h89b, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89a, 12'h789, 12'h99a, 12'habb, 12'h999, 12'h556, 12'h555, 12'h556, 12'h556, 12'h667, 12'h789, 12'h78a, 12'h789, 12'h78a, 12'h79b, 12'h79b, 12'h79b, 12'h89c, 12'h8ac, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hacd, 12'h8ab, 12'h567, 12'h678, 12'h79b, 12'h9ad, 12'hbcd, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hbce, 12'haad, 12'habd, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'h9ad, 12'h8ac, 12'h89c, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h89c, 12'h9ac, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h99c, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hccc, 12'hdde, 12'hfff, 12'heff, 12'hddd, 12'hccd, 12'hccd, 12'hccd, 12'hbcd, 12'habc, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ab, 12'h99b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h89b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'hbbd, 12'h89a, 12'h88a, 12'h99b, 12'h99b, 12'hbcd, 12'h9ab, 12'habc, 12'hcce, 12'hcce, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 
12'habd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habd, 12'habd, 12'habd, 12'haac, 12'haac, 12'haac, 12'h9ab, 12'h89a, 12'h88a, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h89a, 12'h88a, 12'h789, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h677, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h676, 12'h787, 12'h999, 12'habb, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hddd, 12'hcbb, 12'h888, 12'h888, 12'h888, 12'h777, 12'h556, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h666, 12'h566, 12'h556, 12'h556, 12'h456, 12'h455, 12'h455, 12'h455, 12'h444, 12'h344, 12'h344, 12'h245, 12'h456, 12'h568, 12'h689, 12'h78a, 12'h69a, 12'h79b, 12'h79b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h77a, 12'h67a, 12'h67a, 12'h78b, 12'h89c, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h89b, 12'h57a, 12'h46a, 12'h46a, 12'h57b, 12'h79c, 12'h8ad, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h9be, 12'h8be, 12'h8bf, 12'h8be, 12'h8bf, 12'h8be, 12'h8be, 12'h8be, 
12'h8be, 12'h7ae, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h69c, 12'h69c, 12'h69c, 12'h68c, 12'h68c, 12'h68c, 12'h68c, 12'h68b, 12'h68b, 12'h68b, 12'h67a, 12'h57a, 12'h579, 12'h569, 12'h458, 12'h346, 12'h345, 12'h345, 12'h244, 12'h234, 12'h234, 12'h344, 12'h344, 12'h334, 12'h334, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h446, 12'h556, 12'h667, 12'h788, 12'h99a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccb, 12'h999, 12'h877, 12'h777, 12'h666, 12'h666, 12'h677, 12'h778, 12'h89a, 12'hacd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 
12'h9ab, 12'h89b, 12'h88a, 12'h9ab, 12'hbbc, 12'hccc, 12'hccc, 12'h777, 12'h555, 12'h566, 12'h555, 12'h555, 12'h556, 12'h677, 12'h899, 12'h899, 12'h778, 12'h89b, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h8ac, 12'h8ac, 12'h79a, 12'h789, 12'h88a, 12'h88a, 12'h678, 12'h667, 12'h677, 12'h678, 12'h678, 12'h789, 12'h78a, 12'h79b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'h9ce, 12'h9be, 12'h8ab, 12'h678, 12'h678, 12'h78a, 12'h89c, 12'hcde, 12'heff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'habd, 12'habd, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbcf, 12'hccf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hcdf, 12'hccf, 12'hccf, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcce, 12'hbce, 12'hbce, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'h9ad, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h78b, 12'h78b, 12'h78b, 12'h88b, 12'habc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccc, 12'hdde, 12'hfff, 12'hfff, 12'hddd, 12'hccd, 12'hccd, 12'hccd, 12'hbbc, 12'habc, 12'habc, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'haac, 12'haac, 12'hbbc, 12'h99b, 12'h88a, 12'h89a, 12'haab, 12'hccd, 12'h568, 12'h578, 12'h89a, 12'h99b, 12'hbcd, 12'hcce, 12'habd, 12'hbbd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hace, 12'hace, 12'hace, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h99b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h789, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h677, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hbbc, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hedd, 12'hccc, 12'h999, 12'h888, 12'h888, 12'h777, 12'h556, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h666, 12'h556, 12'h556, 12'h456, 12'h456, 12'h455, 12'h455, 12'h445, 12'h445, 12'h344, 12'h245, 12'h346, 12'h467, 12'h689, 12'h78a, 12'h79a, 12'h79b, 12'h79b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h89b, 12'h78a, 12'h77a, 12'h67a, 12'h78b, 12'h78b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h78b, 12'h57a, 12'h46a, 12'h46b, 12'h68c, 12'h79d, 12'h8ae, 12'h8be, 12'h8be, 12'h9be, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h8be, 12'h8be, 
12'h8be, 12'h7be, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h79d, 12'h69c, 12'h69c, 12'h69c, 12'h69c, 12'h68c, 12'h68c, 12'h68c, 12'h68c, 12'h78c, 12'h78b, 12'h68b, 12'h67a, 12'h67a, 12'h679, 12'h568, 12'h457, 12'h346, 12'h235, 12'h234, 12'h234, 12'h234, 12'h344, 12'h344, 12'h334, 12'h344, 12'h445, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h778, 12'h889, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h777, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h899, 12'hacd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcef, 12'hcdf, 12'hcef, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbcd, 
12'hbbd, 12'habd, 12'haac, 12'h89b, 12'h89b, 12'haab, 12'hbbc, 12'h99a, 12'h666, 12'h566, 12'h566, 12'h566, 12'h666, 12'h778, 12'h889, 12'h889, 12'h789, 12'h9ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h89b, 12'h79b, 12'h89b, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'h9ce, 12'h9ce, 12'hace, 12'h9ce, 12'h9bd, 12'h8ab, 12'h678, 12'h678, 12'h78a, 12'h8ac, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hcdd, 12'hbbd, 12'hbbe, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hbce, 12'hccf, 12'hcdf, 12'hccf, 12'hccf, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'haad, 12'h9ad, 12'h89c, 12'h79b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ad, 
12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h78b, 12'h78b, 12'h78b, 12'h89c, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hddd, 12'hccd, 12'hccd, 12'hbbd, 12'habc, 12'habc, 12'habd, 12'habd, 12'h9bd, 12'haad, 12'haad, 12'haad, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haad, 12'haad, 12'habd, 12'haac, 12'h78a, 12'h88a, 12'haac, 12'haac, 12'habc, 12'h679, 12'h457, 12'h457, 12'h568, 12'hdde, 12'hdde, 12'hbcd, 12'hdde, 12'hccd, 12'h89a, 12'h88a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89a, 12'h89b, 
12'h89b, 12'h99b, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ab, 12'h89b, 12'h88a, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h789, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h666, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h888, 12'h888, 12'h777, 12'h666, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h666, 12'h556, 12'h556, 12'h456, 12'h456, 12'h556, 12'h455, 12'h445, 12'h445, 12'h345, 12'h345, 12'h245, 12'h357, 12'h578, 12'h68a, 12'h79a, 12'h79b, 12'h8ab, 12'h8ab, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h89c, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h68a, 12'h57a, 12'h47b, 12'h47b, 12'h79d, 12'h8ae, 12'h8be, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h8be, 
12'h8be, 12'h8be, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h79c, 12'h79c, 12'h79c, 12'h69c, 12'h69c, 12'h79c, 12'h79c, 12'h69c, 12'h68c, 12'h68b, 12'h68b, 12'h68b, 12'h67a, 12'h67a, 12'h679, 12'h457, 12'h446, 12'h445, 12'h335, 12'h334, 12'h334, 12'h344, 12'h334, 12'h334, 12'h334, 12'h345, 12'h456, 12'h556, 12'h567, 12'h668, 12'h779, 12'h789, 12'h779, 12'h668, 12'h668, 12'h788, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'ha99, 12'h888, 12'h889, 12'h778, 12'h667, 12'h777, 12'h777, 12'h899, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 12'hbce, 
12'hbce, 12'hbcd, 12'habd, 12'h9ac, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h788, 12'h778, 12'h778, 12'h789, 12'h789, 12'h78a, 12'h89a, 12'h8ab, 12'h9ac, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'h9ce, 12'hace, 12'hace, 12'h9ce, 12'h9bd, 12'h8ab, 12'h677, 12'h678, 12'h78b, 12'h9bd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hccf, 12'hcdf, 12'hccf, 12'hbcf, 12'hbcf, 12'hbcf, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hbce, 12'hbce, 12'hbcf, 12'hbce, 12'hccf, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'h9ad, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ad, 12'habd, 
12'habd, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h89b, 12'h78b, 12'h77b, 12'h9ac, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'heee, 12'hfff, 12'heff, 12'hddd, 12'hccd, 12'hccd, 12'hbbc, 12'habc, 12'habc, 12'haad, 12'haad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'h99b, 12'h88a, 12'haac, 12'haad, 12'habd, 12'hbbd, 12'hbcd, 12'haac, 12'h678, 12'h789, 12'hbbc, 12'hbbc, 12'hbcd, 12'hccd, 12'hbbd, 12'h9ab, 12'h89a, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h789, 12'h779, 12'h779, 
12'h779, 12'h779, 12'h78a, 12'h89b, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h99b, 12'h89a, 12'h88a, 12'h78a, 12'h77a, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h88a, 12'h789, 12'h778, 12'h778, 12'h677, 12'h677, 12'h777, 12'h777, 12'h777, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h665, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hbbb, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h888, 12'h778, 12'h666, 12'h555, 12'h445, 12'h445, 12'h445, 12'h345, 12'h445, 12'h455, 12'h556, 12'h556, 12'h556, 12'h456, 12'h556, 12'h556, 12'h455, 12'h445, 12'h445, 12'h344, 12'h345, 12'h345, 12'h456, 12'h567, 12'h678, 12'h789, 12'h79a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ab, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h78a, 12'h78a, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h89c, 12'h89c, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h68b, 12'h57a, 12'h47a, 12'h47b, 12'h58c, 12'h7ad, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 
12'h8be, 12'h8bd, 12'h8ad, 12'h7ad, 12'h7ad, 12'h7ac, 12'h7ad, 12'h7ac, 12'h7ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h69c, 12'h69c, 12'h68b, 12'h68b, 12'h68a, 12'h67a, 12'h679, 12'h558, 12'h446, 12'h446, 12'h335, 12'h334, 12'h334, 12'h334, 12'h334, 12'h234, 12'h234, 12'h334, 12'h345, 12'h456, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h88a, 12'h779, 12'h667, 12'h778, 12'h99a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbcd, 12'hbce, 12'h9ac, 12'h788, 12'h777, 12'h778, 12'h899, 12'habc, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hbce, 
12'hbce, 12'hbce, 12'hbcd, 12'habd, 12'h9bc, 12'h9ac, 12'h9ab, 12'h89b, 12'h89b, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'hacd, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'h9cd, 12'h9bd, 12'h8ab, 12'h667, 12'h679, 12'h79b, 12'habd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hccf, 12'hbcf, 12'hbcf, 12'hccf, 12'hccf, 12'hbcf, 12'hccf, 12'hccf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h99c, 12'h78b, 12'h78b, 12'hbbd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdee, 12'hccc, 12'hccd, 12'hfff, 12'hfff, 12'hddd, 12'hccd, 12'hbbc, 12'habc, 12'habc, 12'haac, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'haac, 12'h89a, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h9ac, 12'hbce, 12'hcce, 12'habc, 12'habc, 12'haab, 12'hbcd, 12'hcde, 12'hcce, 12'hbcd, 12'hbcd, 12'habd, 12'haac, 12'h99b, 12'h78a, 12'h779, 12'h789, 12'h889, 12'h889, 12'h789, 
12'h779, 12'h678, 12'h568, 12'h568, 12'h678, 12'h78a, 12'h9ab, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'haad, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88a, 12'h88a, 12'h78a, 12'h78a, 12'h89b, 12'h99c, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h89a, 12'h789, 12'h778, 12'h778, 12'h677, 12'h667, 12'h677, 12'h777, 12'h777, 12'h677, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h666, 12'h766, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'h888, 12'h888, 12'h888, 12'h777, 12'h556, 12'h455, 12'h445, 12'h345, 12'h345, 12'h445, 12'h445, 12'h556, 12'h556, 12'h455, 12'h456, 12'h456, 12'h556, 12'h455, 12'h445, 12'h345, 12'h344, 12'h335, 12'h345, 12'h356, 12'h456, 12'h467, 12'h578, 12'h679, 12'h689, 12'h689, 12'h68a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h68a, 12'h67a, 12'h67a, 12'h67a, 12'h68a, 12'h78b, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h79b, 12'h58b, 12'h47a, 12'h47b, 12'h58b, 12'h79d, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9be, 12'h8be, 12'h8be, 12'h8bd, 
12'h8bd, 12'h8bd, 12'h8ac, 12'h8ac, 12'h7ac, 12'h7ac, 12'h7ac, 12'h7ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h69b, 12'h68b, 12'h67a, 12'h679, 12'h568, 12'h457, 12'h446, 12'h446, 12'h335, 12'h334, 12'h335, 12'h335, 12'h334, 12'h334, 12'h234, 12'h234, 12'h234, 12'h345, 12'h346, 12'h456, 12'h567, 12'h789, 12'h88a, 12'h889, 12'h667, 12'h778, 12'h889, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hcde, 12'hdef, 12'hddf, 12'hbce, 12'h89a, 12'h777, 12'h777, 12'h889, 12'habc, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hcde, 12'hcde, 
12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h9ce, 12'h8ab, 12'h567, 12'h689, 12'h89c, 12'habd, 12'hdde, 12'heff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hcce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hccf, 12'hbcf, 12'hccf, 12'hccf, 12'hbcf, 12'hbcf, 12'hbcf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'haad, 12'h89c, 12'h9ac, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hcdd, 12'haab, 12'hccc, 12'heef, 12'hdde, 12'hccd, 12'hbbc, 12'hbbc, 12'habc, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haac, 12'haac, 12'h9ab, 12'h88a, 12'h88a, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'haac, 12'hccd, 12'hccd, 12'haac, 12'hbcd, 12'hcce, 12'hcce, 12'hbcd, 12'hbbd, 12'habc, 12'haac, 12'h9ac, 12'h88a, 12'h779, 12'h779, 12'h88a, 12'h99a, 12'h99a, 
12'h99a, 12'h899, 12'h889, 12'h778, 12'h667, 12'h457, 12'h568, 12'h78a, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'haad, 12'haac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89b, 12'h99b, 12'h99b, 12'h89a, 12'h789, 12'h778, 12'h778, 12'h677, 12'h667, 12'h677, 12'h777, 12'h777, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h555, 12'h555, 12'h655, 12'h555, 12'h555, 12'h655, 12'h665, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hbbb, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h888, 12'h778, 12'h777, 12'h566, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h334, 12'h334, 12'h334, 12'h344, 12'h245, 12'h356, 12'h356, 12'h356, 12'h467, 12'h568, 12'h568, 12'h578, 12'h679, 12'h679, 12'h679, 12'h67a, 12'h68a, 12'h679, 12'h579, 12'h579, 12'h68a, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h79b, 12'h68b, 12'h57a, 12'h47b, 12'h57b, 12'h69c, 12'h8ad, 12'h9be, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9ce, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bc, 
12'h8ac, 12'h8ac, 12'h7ac, 12'h7ac, 12'h7ac, 12'h79c, 12'h7ac, 12'h7ac, 12'h79c, 12'h69b, 12'h69b, 12'h69b, 12'h79c, 12'h7ac, 12'h79c, 12'h79b, 12'h69b, 12'h68a, 12'h67a, 12'h679, 12'h669, 12'h568, 12'h447, 12'h447, 12'h346, 12'h345, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h234, 12'h234, 12'h345, 12'h345, 12'h346, 12'h446, 12'h567, 12'h779, 12'h899, 12'h778, 12'h678, 12'h889, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdef, 12'hcdf, 12'hcdf, 12'hbde, 12'h9ab, 12'h788, 12'h677, 12'h788, 12'haac, 12'hbde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hcdf, 12'hcde, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h9bd, 12'h8ab, 12'h677, 12'h689, 12'h9bd, 12'hacd, 12'hdde, 12'heff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbce, 12'hbce, 12'hccf, 12'hbce, 12'hbce, 12'hbcf, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ad, 12'h99c, 12'haad, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccc, 12'h99a, 12'haab, 12'hccc, 12'hccd, 12'hbbc, 12'hbbc, 12'habc, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haac, 12'haac, 12'h99b, 12'h78a, 12'h679, 12'h89b, 12'h9ac, 12'h9ad, 12'habe, 12'hbbe, 12'habd, 12'h99c, 12'h88b, 12'haac, 12'h99b, 12'habc, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'h9ac, 12'h9ac, 12'h99b, 12'h88a, 12'h88a, 12'h99a, 12'haab, 12'haab, 
12'h99a, 12'h788, 12'h888, 12'h899, 12'h899, 12'h788, 12'h778, 12'h689, 12'h679, 12'h78a, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h99b, 12'h99b, 12'h99b, 12'h889, 12'h778, 12'h778, 12'h677, 12'h677, 12'h677, 12'h777, 12'h777, 12'h677, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h656, 12'h556, 12'h655, 12'h655, 12'h655, 12'h655, 12'h665, 12'h666, 12'h776, 12'h887, 12'h999, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h888, 12'h777, 12'h677, 12'h556, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h344, 12'h344, 12'h334, 12'h234, 12'h244, 12'h245, 12'h355, 12'h355, 12'h456, 12'h456, 12'h457, 12'h567, 12'h678, 12'h679, 12'h689, 12'h679, 12'h679, 12'h579, 12'h67a, 12'h57a, 12'h68a, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h68b, 12'h57a, 12'h57b, 12'h58b, 12'h68c, 12'h8ad, 12'h9be, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9ce, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bc, 12'h8ac, 12'h8ab, 
12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h89b, 12'h89b, 12'h79b, 12'h78b, 12'h68a, 12'h68b, 12'h79b, 12'h79b, 12'h79b, 12'h68a, 12'h579, 12'h569, 12'h569, 12'h669, 12'h669, 12'h669, 12'h558, 12'h558, 12'h457, 12'h346, 12'h346, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h234, 12'h345, 12'h346, 12'h346, 12'h346, 12'h456, 12'h667, 12'h889, 12'h778, 12'h778, 12'h889, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcde, 12'habe, 12'h9ad, 12'h9bd, 12'h89b, 12'h788, 12'h677, 12'h788, 12'h9ab, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hcde, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h9bd, 12'h8ab, 12'h677, 12'h78a, 12'hace, 12'hbce, 12'hdde, 12'heff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hcdf, 12'hddf, 12'hcdf, 12'hccf, 12'hcdf, 12'hccf, 12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbcf, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbbe, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ad, 12'h9ac, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbbc, 12'haab, 12'h99a, 12'haab, 12'hbbc, 12'hbbc, 12'habc, 12'habc, 12'haad, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h88a, 12'h568, 12'h78a, 12'h9ac, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'h99c, 12'h9ac, 12'h78a, 12'haac, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h99b, 12'h9ab, 12'haab, 
12'h889, 12'h566, 12'h566, 12'h787, 12'h999, 12'h999, 12'h99a, 12'h9aa, 12'h99a, 12'h88a, 12'h78a, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h99b, 12'h89b, 12'h88a, 12'h779, 12'h778, 12'h777, 12'h677, 12'h677, 12'h777, 12'h777, 12'h777, 12'h677, 12'h677, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h655, 12'h655, 12'h655, 12'h665, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h677, 12'h566, 12'h555, 12'h445, 12'h445, 12'h445, 12'h345, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h344, 12'h334, 12'h344, 12'h344, 12'h344, 12'h345, 12'h345, 12'h456, 12'h456, 12'h457, 12'h567, 12'h578, 12'h679, 12'h789, 12'h678, 12'h568, 12'h568, 12'h67a, 12'h68a, 12'h78b, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h79b, 12'h79b, 12'h68b, 12'h68b, 12'h68b, 12'h79c, 12'h8ad, 12'h9be, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9ce, 12'h9cd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bc, 12'h8ac, 12'h8ab, 12'h89b, 12'h79a, 
12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79a, 12'h78a, 12'h79a, 12'h79a, 12'h78a, 12'h579, 12'h458, 12'h458, 12'h558, 12'h569, 12'h66a, 12'h669, 12'h569, 12'h569, 12'h568, 12'h457, 12'h456, 12'h456, 12'h445, 12'h335, 12'h334, 12'h334, 12'h345, 12'h345, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h557, 12'h778, 12'h778, 12'h778, 12'h888, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hcde, 12'h8ad, 12'h78c, 12'h89c, 12'h9ac, 12'h899, 12'h778, 12'h788, 12'h9ab, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcde, 
12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h9bd, 12'h8ac, 12'h678, 12'h79a, 12'h9be, 12'hbce, 12'hdde, 12'heff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hcdf, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbcf, 12'hbcf, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ad, 12'haad, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbcc, 12'hbbc, 12'haab, 12'h99b, 12'h99a, 12'h9ab, 12'haac, 12'habc, 12'habc, 12'haac, 12'haac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'h89b, 12'h679, 12'h78a, 12'h9ac, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'h9ac, 12'haac, 12'h89a, 12'h89a, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbce, 12'hbce, 12'hbbd, 12'haac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 
12'h89a, 12'h778, 12'h666, 12'h676, 12'h787, 12'h898, 12'h999, 12'h999, 12'h9aa, 12'haab, 12'habc, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h99c, 12'h9ac, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h88a, 12'h779, 12'h778, 12'h677, 12'h677, 12'h677, 12'h777, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h655, 12'h665, 12'h666, 12'h766, 12'h777, 12'h888, 12'haaa, 12'hbbc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccb, 12'h888, 12'h666, 12'h555, 12'h455, 12'h445, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h344, 12'h444, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h444, 12'h344, 12'h344, 12'h334, 12'h345, 12'h345, 12'h445, 12'h446, 12'h456, 12'h567, 12'h567, 12'h678, 12'h679, 12'h568, 12'h457, 12'h458, 12'h579, 12'h67a, 12'h78b, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h78b, 12'h68b, 12'h78b, 12'h79c, 12'h89d, 12'h9ad, 12'h9bd, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bc, 12'h9bc, 12'h8ab, 12'h8ab, 12'h89a, 12'h789, 12'h789, 12'h779, 
12'h779, 12'h779, 12'h78a, 12'h88a, 12'h89b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h79a, 12'h78a, 12'h78a, 12'h67a, 12'h569, 12'h458, 12'h459, 12'h569, 12'h66a, 12'h67b, 12'h67b, 12'h77b, 12'h78a, 12'h67a, 12'h568, 12'h557, 12'h447, 12'h446, 12'h345, 12'h335, 12'h345, 12'h345, 12'h345, 12'h346, 12'h446, 12'h446, 12'h346, 12'h346, 12'h456, 12'h668, 12'h778, 12'h678, 12'h888, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hcde, 12'h8ae, 12'h79d, 12'hbce, 12'hbde, 12'h9ab, 12'h788, 12'h788, 12'h9ab, 12'hbcd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcde, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h9bd, 12'h8ab, 12'h678, 12'h78a, 12'h9bd, 12'hace, 12'hdde, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'haad, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hcdf, 12'hddf, 12'hcdf, 12'hccf, 12'hccf, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbcf, 12'hbcf, 12'hbcf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ad, 12'hbbd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcc, 12'habc, 12'habc, 12'habc, 12'h9ab, 12'h89a, 12'h89a, 12'h89a, 12'h9ab, 12'haac, 12'haac, 12'haac, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'h9ac, 12'h679, 12'h78a, 12'haad, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'h99b, 12'h88a, 12'h99a, 12'haac, 12'hbbd, 12'hbbd, 12'hbce, 12'hcce, 12'hbce, 12'habd, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h9ab, 12'haac, 12'haac, 
12'haab, 12'h99b, 12'h89a, 12'h889, 12'h788, 12'h787, 12'h898, 12'h898, 12'h888, 12'h788, 12'h99a, 12'haab, 12'hbbc, 12'hbbc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h88a, 12'h778, 12'h678, 12'h677, 12'h677, 12'h677, 12'h777, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h566, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h334, 12'h334, 12'h445, 12'h445, 12'h456, 12'h456, 12'h456, 12'h557, 12'h567, 12'h678, 12'h678, 12'h568, 12'h458, 12'h348, 12'h459, 12'h67a, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h68b, 12'h68b, 12'h78b, 12'h78c, 12'h89c, 12'h89c, 12'h9ad, 12'h9ad, 12'habe, 12'habe, 12'habe, 12'hace, 12'hace, 12'hace, 12'hace, 12'hacd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bc, 12'h9ab, 12'h8ab, 12'h79a, 12'h789, 12'h779, 12'h778, 12'h769, 12'h879, 
12'h88a, 12'h99a, 12'haab, 12'haab, 12'habc, 12'habb, 12'haab, 12'h9ab, 12'h9ab, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h67a, 12'h569, 12'h569, 12'h67a, 12'h67b, 12'h78c, 12'h78c, 12'h78c, 12'h78b, 12'h78b, 12'h78b, 12'h67a, 12'h568, 12'h447, 12'h447, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h456, 12'h457, 12'h457, 12'h446, 12'h246, 12'h456, 12'h668, 12'h678, 12'h678, 12'h788, 12'h9aa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hdde, 12'h9ae, 12'h8ad, 12'hcdf, 12'hdef, 12'hacd, 12'h789, 12'h778, 12'h89a, 12'hacd, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hcde, 
12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'hace, 12'h9ce, 12'h9bd, 12'h9bd, 12'h89b, 12'h678, 12'h79b, 12'h8ad, 12'h9bd, 12'hcde, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'habe, 12'hbce, 12'hcce, 12'hccf, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hccf, 12'hccf, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbbe, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ad, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbcd, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h89b, 12'h88a, 12'h89b, 12'h9ab, 12'haac, 12'habc, 12'habd, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'haac, 12'haac, 12'h78a, 12'h77a, 12'haac, 12'hbbe, 12'hbce, 12'hccf, 12'hccf, 12'hbce, 12'habe, 12'habe, 12'habd, 12'haad, 12'haad, 12'h88b, 12'h88a, 12'h99b, 12'h89b, 12'haac, 12'hbbd, 12'hbbd, 12'hbce, 12'hbce, 12'hbbe, 12'haad, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'haac, 
12'haac, 12'haac, 12'haac, 12'haab, 12'h99a, 12'h89a, 12'h899, 12'h899, 12'h788, 12'h677, 12'h667, 12'h789, 12'h89a, 12'h89a, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89a, 12'h779, 12'h678, 12'h677, 12'h677, 12'h677, 12'h777, 12'h777, 12'h667, 12'h677, 12'h667, 12'h666, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hddc, 12'h999, 12'h666, 12'h555, 12'h455, 12'h455, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h334, 12'h335, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h467, 12'h568, 12'h678, 12'h679, 12'h679, 12'h669, 12'h569, 12'h459, 12'h569, 12'h78b, 12'h89b, 12'h89c, 12'h79b, 12'h78b, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h99d, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'hace, 12'hacd, 12'hacd, 12'hacd, 12'h9bd, 12'h9bd, 12'h9bc, 12'h9bc, 12'h8ab, 12'h89a, 12'h789, 12'h678, 12'h678, 12'h779, 12'h879, 12'h88a, 12'h99b, 
12'haab, 12'hbbc, 12'hbbc, 12'hbbc, 12'habc, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h8ab, 12'h8ab, 12'h89b, 12'h89b, 12'h79b, 12'h67a, 12'h56a, 12'h57a, 12'h78b, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h78c, 12'h78b, 12'h78b, 12'h68a, 12'h569, 12'h358, 12'h357, 12'h357, 12'h346, 12'h346, 12'h346, 12'h456, 12'h557, 12'h567, 12'h567, 12'h457, 12'h346, 12'h457, 12'h668, 12'h678, 12'h678, 12'h778, 12'h99a, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdef, 12'h9be, 12'habe, 12'hdef, 12'hdef, 12'hcdf, 12'h9ab, 12'h778, 12'h889, 12'habc, 12'hbde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'heef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hcde, 
12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hcdf, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hbcf, 12'habe, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h89b, 12'h689, 12'h89b, 12'h8ac, 12'h9bd, 12'hbce, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h9ad, 12'habd, 12'hbce, 12'hbce, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'haad, 12'h9ac, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'h89b, 12'h77a, 12'h9ac, 12'hbbd, 12'hbbe, 12'hccf, 12'hccf, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'haad, 12'haad, 12'h78a, 12'h88a, 12'h88a, 12'h779, 12'h9ac, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbd, 12'habd, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h88b, 12'h89b, 
12'h99b, 12'haac, 12'haac, 12'habc, 12'habc, 12'h9ab, 12'h99a, 12'h89a, 12'h899, 12'h788, 12'h678, 12'h678, 12'h789, 12'h88a, 12'h88a, 12'h789, 12'h88a, 12'h99b, 12'h9ac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h89a, 12'h789, 12'h678, 12'h677, 12'h677, 12'h777, 12'h777, 12'h777, 12'h667, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h665, 12'h666, 12'h766, 12'h777, 12'h988, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h777, 12'h566, 12'h455, 12'h455, 12'h445, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h335, 12'h335, 12'h345, 12'h445, 12'h446, 12'h456, 12'h557, 12'h567, 12'h678, 12'h679, 12'h78a, 12'h78a, 12'h78b, 12'h78b, 12'h67a, 12'h569, 12'h78b, 12'h9ac, 12'h9ad, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bc, 12'h9bc, 12'h8ab, 12'h79a, 12'h789, 12'h689, 12'h678, 12'h778, 12'h889, 12'h99a, 12'h99a, 12'haab, 12'hbbc, 
12'hbbc, 12'hccc, 12'hbcc, 12'hbbc, 12'haab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h8ab, 12'h8ab, 12'h8ab, 12'h89b, 12'h89b, 12'h79b, 12'h68b, 12'h57a, 12'h68b, 12'h79c, 12'h8ad, 12'h89d, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h69b, 12'h57a, 12'h369, 12'h258, 12'h357, 12'h357, 12'h346, 12'h346, 12'h457, 12'h568, 12'h678, 12'h678, 12'h567, 12'h356, 12'h457, 12'h678, 12'h778, 12'h778, 12'h778, 12'h999, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'habe, 12'hbcf, 12'hdef, 12'hcdf, 12'hcdf, 12'habd, 12'h788, 12'h789, 12'habc, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hcdf, 12'hcde, 
12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hcce, 12'hcdf, 12'hddf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hace, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h89b, 12'h68a, 12'h8ac, 12'h8ac, 12'h9ad, 12'hbce, 12'hdde, 12'heff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'h9ad, 12'h89c, 12'h78b, 12'h89c, 12'h9ad, 12'habd, 12'hbce, 12'hbce, 12'hccf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbbe, 12'haad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h9ad, 12'h9ad, 12'habd, 12'hbce, 12'hbce, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'haac, 12'habd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccd, 12'hbbc, 12'haac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h88a, 12'h78a, 12'h88a, 12'h89b, 12'h89b, 12'h88b, 12'h88a, 12'h9ac, 12'hbbd, 12'hbbd, 12'hbce, 12'hcdf, 12'hbcf, 12'habe, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h78a, 12'h78a, 12'h88a, 12'h78a, 12'h99b, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h78a, 
12'h78a, 12'h89b, 12'h89b, 12'h9ac, 12'haac, 12'haac, 12'h9ab, 12'h9ab, 12'h9ab, 12'h89a, 12'h789, 12'h789, 12'h779, 12'h789, 12'h89a, 12'h678, 12'h557, 12'h789, 12'h99a, 12'h9ab, 12'haab, 12'haac, 12'haac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89b, 12'h99b, 12'h89a, 12'h889, 12'h778, 12'h677, 12'h778, 12'h778, 12'h777, 12'h777, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h665, 12'h666, 12'h666, 12'h777, 12'h888, 12'h999, 12'haaa, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'h999, 12'h666, 12'h455, 12'h445, 12'h445, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h444, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h334, 12'h345, 12'h345, 12'h345, 12'h456, 12'h556, 12'h567, 12'h568, 12'h679, 12'h78a, 12'h78a, 12'h78b, 12'h89b, 12'h89c, 12'h89b, 12'h68a, 12'h79b, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h8ab, 12'h79a, 12'h689, 12'h678, 12'h678, 12'h778, 12'h889, 12'h9aa, 12'habb, 12'habb, 12'hbbc, 12'hbbc, 
12'hbcc, 12'hccc, 12'hbbc, 12'haab, 12'h9ab, 12'h9ab, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h68b, 12'h57a, 12'h68b, 12'h79c, 12'h8ad, 12'h89d, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h58b, 12'h47a, 12'h258, 12'h358, 12'h357, 12'h457, 12'h457, 12'h457, 12'h568, 12'h679, 12'h779, 12'h668, 12'h457, 12'h457, 12'h678, 12'h778, 12'h778, 12'h778, 12'h999, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hbce, 12'hddf, 12'hdef, 12'hddf, 12'hbce, 12'habe, 12'h89a, 12'h788, 12'h9ab, 12'hbce, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcde, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hace, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h89b, 12'h79b, 12'h8ac, 12'h8ac, 12'h9ad, 12'hbce, 12'hdde, 12'heef, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h89c, 12'h78b, 12'h89c, 12'habd, 12'hbbe, 12'hbce, 12'hcce, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hbce, 12'hccf, 12'hccf, 12'hbce, 12'hbce, 12'hbbe, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ad, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdde, 12'hccd, 12'hbbc, 12'haac, 12'h9ac, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88b, 12'h78a, 12'h88b, 12'h9ac, 12'habd, 12'habd, 12'hbbe, 12'hccf, 12'hcdf, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h89b, 12'h779, 12'h99b, 12'h99b, 12'h99c, 12'h9ac, 12'habd, 12'habd, 12'hbbd, 12'hbbe, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h99b, 
12'h88b, 12'h78a, 12'h78b, 12'h78b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h89b, 12'h89a, 12'h88a, 12'h88a, 12'h89a, 12'h778, 12'h567, 12'h889, 12'h899, 12'h89a, 12'h89a, 12'h89a, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h99b, 12'h89a, 12'h889, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h667, 12'h667, 12'h677, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h777, 12'h555, 12'h444, 12'h445, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h457, 12'h468, 12'h468, 12'h569, 12'h78a, 12'h78b, 12'h89b, 12'h89c, 12'h9ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h89a, 12'h789, 12'h678, 12'h678, 12'h789, 12'h89a, 12'h9ab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 
12'hbbc, 12'hbbc, 12'habb, 12'h9aa, 12'h99a, 12'h89a, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h79b, 12'h79b, 12'h78b, 12'h68b, 12'h57b, 12'h68b, 12'h79c, 12'h8ad, 12'h79d, 12'h79c, 12'h79c, 12'h79c, 12'h79d, 12'h7ad, 12'h79c, 12'h68c, 12'h57a, 12'h469, 12'h358, 12'h358, 12'h457, 12'h457, 12'h457, 12'h568, 12'h679, 12'h679, 12'h568, 12'h457, 12'h457, 12'h668, 12'h678, 12'h668, 12'h778, 12'h999, 12'hbbc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hcdf, 12'hdef, 12'hdef, 12'hbcf, 12'h9ad, 12'h8ad, 12'h9ab, 12'h789, 12'h9ab, 12'hbce, 12'hcde, 12'hbde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hcde, 12'hcde, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hbce, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ac, 12'h9ad, 12'hbce, 12'hdee, 12'heff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h99c, 12'h78b, 12'h78b, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habd, 12'h9ad, 12'h9ad, 12'h89c, 12'h78b, 12'h89c, 12'h9ac, 12'habd, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'hbcd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h78b, 12'h88b, 12'h78b, 12'h78b, 12'h89b, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hcdf, 12'hccf, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h99b, 12'h78a, 12'h99b, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haac, 
12'h9ac, 12'h99c, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ac, 12'h9ab, 12'h89b, 12'h99b, 12'h99b, 12'h678, 12'h668, 12'h889, 12'h899, 12'h89a, 12'h899, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h889, 12'h789, 12'h778, 12'h778, 12'h778, 12'h778, 12'h677, 12'h667, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h888, 12'h999, 12'haaa, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h788, 12'h555, 12'h555, 12'h444, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h345, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h457, 12'h568, 12'h568, 12'h569, 12'h568, 12'h569, 12'h78a, 12'h89b, 12'h89b, 12'h89c, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bc, 12'h9bc, 12'h9ac, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h789, 12'h789, 12'h789, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h99a, 12'h99a, 
12'haab, 12'haab, 12'h99a, 12'h88a, 12'h88a, 12'h78a, 12'h78a, 12'h779, 12'h679, 12'h67a, 12'h67a, 12'h68b, 12'h68b, 12'h78b, 12'h68b, 12'h67b, 12'h57b, 12'h79c, 12'h8ad, 12'h8ad, 12'h79c, 12'h79d, 12'h79d, 12'h7ad, 12'h8ad, 12'h79d, 12'h79c, 12'h68b, 12'h56a, 12'h459, 12'h358, 12'h457, 12'h457, 12'h457, 12'h568, 12'h679, 12'h679, 12'h668, 12'h568, 12'h567, 12'h567, 12'h668, 12'h667, 12'h778, 12'h999, 12'hbcc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdef, 12'hcdf, 12'hbce, 12'h9ad, 12'h79c, 12'h89c, 12'h9ac, 12'h899, 12'h89a, 12'hbce, 12'hcdf, 12'hbce, 12'hbde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'hcdf, 12'hcde, 12'hcde, 12'hcce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ac, 12'h9bd, 12'h8ad, 12'h89c, 12'h8ac, 12'hbce, 12'hdee, 12'heff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h89c, 12'h78b, 12'h89c, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h78b, 12'h89c, 12'h9ac, 12'haad, 12'habd, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'hbcd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcd, 12'hbbd, 12'habd, 12'haad, 12'haac, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h88b, 12'h78a, 12'h78a, 12'h78a, 12'h67a, 12'h78a, 12'h78b, 12'h88b, 12'h99c, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hccf, 12'hccf, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h89b, 12'h779, 12'h99b, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'habc, 12'h89b, 12'h557, 12'h779, 12'h88a, 12'h89a, 12'h899, 12'h9ab, 12'hdde, 12'hccd, 12'haab, 12'h89a, 12'h88a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89a, 12'h88a, 12'h889, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h888, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedd, 12'hccc, 12'h888, 12'h666, 12'h555, 12'h444, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h335, 12'h345, 12'h346, 12'h457, 12'h568, 12'h679, 12'h679, 12'h78a, 12'h67a, 12'h579, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bc, 12'h9bc, 12'habd, 12'habc, 12'habd, 12'habd, 12'habc, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9ac, 12'h89b, 12'h79a, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h789, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h98a, 
12'h99b, 12'haab, 12'h88a, 12'h779, 12'h77a, 12'h89a, 12'h88a, 12'h78a, 12'h679, 12'h579, 12'h57a, 12'h57a, 12'h68b, 12'h78b, 12'h78b, 12'h68b, 12'h57b, 12'h79c, 12'h79d, 12'h7ad, 12'h79d, 12'h7ad, 12'h7ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h79d, 12'h78c, 12'h57a, 12'h469, 12'h458, 12'h458, 12'h458, 12'h558, 12'h568, 12'h679, 12'h779, 12'h779, 12'h678, 12'h668, 12'h668, 12'h567, 12'h567, 12'h667, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdef, 12'hbcf, 12'h9ad, 12'h8ad, 12'h89c, 12'h9ad, 12'habd, 12'h9ab, 12'h89a, 12'hbcd, 12'hbde, 12'hbce, 12'hbde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hcde, 12'hcce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ac, 12'h9bd, 12'h8ac, 12'h79c, 12'h89c, 12'habd, 12'hdee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h89c, 12'h78b, 12'h89c, 12'hbbe, 12'hbce, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h88c, 12'h89c, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 
12'hbbe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'hbbd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbcd, 12'habd, 12'haad, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'haac, 12'h9ac, 12'h99b, 12'h89b, 12'h78b, 12'h78a, 12'h67a, 12'h78b, 12'h89c, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hccf, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h99b, 12'h679, 12'h99b, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'haac, 12'habd, 12'habd, 12'habc, 12'hbcd, 12'h89b, 12'h447, 12'h88a, 12'h99b, 12'h89a, 12'h89a, 12'hbbc, 12'hdde, 12'hccd, 12'h899, 12'h667, 12'h668, 12'h778, 12'h88a, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h99b, 12'h99b, 12'h89a, 12'h889, 12'h789, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h677, 12'h667, 12'h667, 12'h677, 12'h677, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h788, 12'h888, 12'haaa, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'hccc, 12'h999, 12'h777, 12'h555, 12'h444, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h345, 12'h445, 12'h445, 12'h445, 12'h346, 12'h346, 12'h447, 12'h558, 12'h679, 12'h78a, 12'h78a, 12'h78b, 12'h78b, 12'h67a, 12'h78b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9ac, 12'h89b, 12'h78a, 12'h78a, 12'h88a, 12'h78a, 12'h88a, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h77a, 12'h88a, 
12'h99b, 12'haac, 12'h88a, 12'h779, 12'h88a, 12'h9ab, 12'h9ab, 12'h99b, 12'h78a, 12'h57a, 12'h56a, 12'h57b, 12'h78b, 12'h78c, 12'h79c, 12'h78c, 12'h57b, 12'h68c, 12'h79d, 12'h7ad, 12'h7ad, 12'h7ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ad, 12'h79c, 12'h68b, 12'h469, 12'h459, 12'h458, 12'h568, 12'h568, 12'h668, 12'h779, 12'h78a, 12'h78a, 12'h68a, 12'h679, 12'h679, 12'h568, 12'h557, 12'h667, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hbce, 12'h9ad, 12'h9ad, 12'h8ac, 12'habd, 12'hcdf, 12'hbcd, 12'h9ab, 12'hbcd, 12'hbce, 12'hbce, 12'hbde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ac, 12'h8ad, 12'h8ad, 12'h79c, 12'h8ac, 12'hbce, 12'hdee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'habd, 12'h9ad, 12'h89c, 12'h89c, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 
12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h88b, 12'h78a, 12'h89b, 12'h9ad, 12'habd, 12'haad, 12'haad, 12'haad, 12'habd, 12'hbbe, 12'hbce, 12'hcce, 12'hbce, 12'habe, 12'habd, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'h9ac, 12'h67a, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'h679, 12'h89a, 12'hbcd, 12'habc, 12'haac, 12'haab, 12'habc, 12'hbbc, 12'haab, 12'h778, 12'h667, 12'h667, 12'h667, 12'h667, 12'h778, 12'h789, 12'h89a, 12'h99b, 12'h99b, 12'h99a, 12'h89a, 12'h889, 12'h788, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h677, 12'h677, 12'h667, 12'h777, 12'h777, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h888, 12'h999, 12'hbbc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h777, 12'h555, 12'h444, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h345, 12'h445, 12'h445, 12'h446, 12'h346, 12'h457, 12'h569, 12'h67a, 12'h78a, 12'h78b, 12'h79b, 12'h89b, 12'h78b, 12'h79b, 12'h89b, 12'h8ac, 12'h9ac, 12'h9ab, 12'h9ac, 12'h8ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h78a, 12'h88a, 12'h89b, 12'h88b, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h87a, 12'h77a, 
12'h98b, 12'haac, 12'h88a, 12'h779, 12'h89a, 12'haac, 12'hbbc, 12'haac, 12'h89b, 12'h68a, 12'h57b, 12'h68b, 12'h79c, 12'h79d, 12'h89d, 12'h89d, 12'h68c, 12'h57b, 12'h79c, 12'h79d, 12'h7ad, 12'h7ae, 12'h8ae, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h7ad, 12'h68b, 12'h46a, 12'h469, 12'h468, 12'h568, 12'h568, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h77a, 12'h568, 12'h457, 12'h667, 12'h99a, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hbce, 12'h9ad, 12'h9ad, 12'h9ad, 12'hbce, 12'hdef, 12'hcde, 12'h9ab, 12'hacd, 12'hbce, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hcdf, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8ac, 12'h7ac, 12'h8ad, 12'h9bd, 12'hace, 12'hcde, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'habd, 12'h9ad, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'haad, 12'h9ad, 12'h9ac, 12'h89c, 12'h9ac, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 
12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hccd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h88b, 12'h99c, 12'habd, 12'haad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hbbe, 12'habd, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'h9ac, 12'h78a, 12'h99b, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'hbce, 12'habc, 12'h89b, 12'hbcd, 12'hbcd, 12'habd, 12'habc, 12'haac, 12'h99a, 12'h889, 12'h778, 12'h778, 12'h677, 12'h667, 12'h677, 12'h667, 12'h667, 12'h667, 12'h678, 12'h778, 12'h889, 12'h889, 12'h889, 12'h788, 12'h788, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h677, 12'h777, 12'h677, 12'h677, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h788, 12'h889, 12'haab, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedd, 12'hbbb, 12'h777, 12'h555, 12'h444, 12'h444, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h445, 12'h344, 12'h345, 12'h345, 12'h446, 12'h447, 12'h458, 12'h579, 12'h68a, 12'h78b, 12'h78b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'h9ab, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h89b, 12'h9ab, 12'h89b, 12'h89a, 12'h89b, 12'h89b, 12'h8ab, 12'h8ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h89a, 12'h89a, 12'h899, 12'h889, 12'h789, 12'h789, 12'h78a, 12'h78a, 12'h79b, 12'h79b, 12'h79b, 12'h89b, 12'h88a, 12'h88b, 12'h99b, 12'haac, 12'h88b, 12'h77a, 
12'h88a, 12'h88a, 12'h779, 12'h779, 12'h99b, 12'habc, 12'habc, 12'h9ac, 12'h89b, 12'h78b, 12'h68c, 12'h79c, 12'h79d, 12'h8ad, 12'h8ae, 12'h8ad, 12'h69c, 12'h47b, 12'h68c, 12'h79d, 12'h7ae, 12'h7ae, 12'h8be, 12'h8be, 12'h8be, 12'h7ae, 12'h7ae, 12'h7ad, 12'h68c, 12'h47a, 12'h469, 12'h468, 12'h568, 12'h568, 12'h679, 12'h78a, 12'h78b, 12'h78b, 12'h89b, 12'h89b, 12'h78a, 12'h568, 12'h457, 12'h668, 12'h99a, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hcdf, 12'h9bd, 12'h9ad, 12'habd, 12'hbce, 12'hdef, 12'hdef, 12'habc, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hbde, 12'hcdf, 12'hcde, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hbcf, 12'hbce, 12'habe, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ac, 12'h79c, 12'h7ac, 12'h9bd, 12'hbde, 12'hcde, 12'heef, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'h9ac, 12'h89c, 12'h89c, 12'h89b, 12'h99c, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbbe, 12'habe, 12'habe, 
12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdde, 12'hccd, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h88b, 12'h89b, 12'haac, 12'haad, 12'h9ad, 12'haad, 12'h9ad, 12'haad, 12'haad, 12'habe, 12'hbbe, 12'hbce, 12'hbce, 12'hbbe, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h88b, 12'h78a, 12'h9ab, 12'habd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 
12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h89b, 12'h9ac, 12'hbcd, 12'habd, 12'haac, 12'h9ac, 12'h99b, 12'h99b, 12'h889, 12'h779, 12'h789, 12'h778, 12'h677, 12'h667, 12'h677, 12'h777, 12'h677, 12'h667, 12'h667, 12'h677, 12'h677, 12'h677, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h888, 12'h999, 12'hccc, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedd, 12'hccc, 12'h888, 12'h555, 12'h444, 12'h444, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h445, 12'h344, 12'h445, 12'h346, 12'h457, 12'h458, 12'h569, 12'h67a, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h78a, 12'h789, 12'h88a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h78a, 12'h789, 12'h78a, 12'h79a, 12'h79a, 12'h79a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h99a, 12'h9aa, 12'h889, 12'h789, 12'h789, 12'h889, 12'h889, 12'h88a, 12'h79a, 12'h78b, 12'h79b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'haac, 12'hbbd, 12'haac, 12'h88a, 
12'h77a, 12'h779, 12'h779, 12'h78a, 12'h9ab, 12'haac, 12'h9ac, 12'h89c, 12'h78b, 12'h78c, 12'h79c, 12'h79d, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h79d, 12'h47b, 12'h58c, 12'h7ad, 12'h7ae, 12'h7be, 12'h8be, 12'h8be, 12'h8be, 12'h7ae, 12'h7ae, 12'h6ad, 12'h69c, 12'h47a, 12'h469, 12'h458, 12'h568, 12'h569, 12'h679, 12'h78b, 12'h78b, 12'h78b, 12'h9ac, 12'h9ac, 12'h89b, 12'h569, 12'h357, 12'h567, 12'h99a, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hcdf, 12'habe, 12'h9ad, 12'h9ad, 12'hbde, 12'hdef, 12'hcef, 12'hbce, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hbde, 12'hcdf, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hcce, 12'hcdf, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ac, 12'h79c, 12'h8ad, 12'hace, 12'hbde, 12'hdde, 12'heff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h99c, 12'h9ac, 12'habd, 12'habd, 12'haad, 12'h78b, 12'h78b, 12'h67a, 12'h68b, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h78b, 12'h78b, 12'h89c, 12'h89c, 12'h89b, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccd, 12'habc, 12'haac, 12'h9ac, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h78a, 12'h77a, 12'h88b, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 
12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'habc, 12'h89b, 12'h9ac, 12'hbbd, 12'habd, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h88a, 12'h889, 12'h778, 12'h678, 12'h677, 12'h667, 12'h666, 12'h677, 12'h667, 12'h667, 12'h666, 12'h667, 12'h667, 12'h677, 12'h777, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h778, 12'h888, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdcc, 12'h999, 12'h666, 12'h444, 12'h444, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h334, 12'h334, 12'h334, 12'h335, 12'h345, 12'h345, 12'h446, 12'h457, 12'h557, 12'h568, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h67a, 12'h78a, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h678, 12'h778, 12'h779, 12'h789, 12'h789, 12'h789, 12'h79a, 12'h789, 12'h789, 12'h789, 12'h778, 12'h678, 12'h678, 12'h778, 12'h889, 12'h889, 12'h788, 12'h778, 12'h788, 12'h789, 12'h88a, 12'h88a, 12'h79b, 12'h78b, 12'h79b, 12'h89b, 12'h9ac, 12'h89b, 12'h89b, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'h99b, 
12'h78a, 12'h77a, 12'h88b, 12'h89b, 12'h99c, 12'h99c, 12'h89c, 12'h89c, 12'h79c, 12'h79d, 12'h79d, 12'h7ad, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 12'h7ad, 12'h48c, 12'h48c, 12'h6ad, 12'h7be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h7be, 12'h7ae, 12'h6ad, 12'h59c, 12'h58b, 12'h369, 12'h459, 12'h458, 12'h469, 12'h57a, 12'h68b, 12'h78b, 12'h78b, 12'h9ac, 12'h9ad, 12'h89c, 12'h569, 12'h357, 12'h668, 12'haaa, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddf, 12'habe, 12'h8ad, 12'h89d, 12'hcdf, 12'hdef, 12'hcdf, 12'hbce, 12'hacd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hace, 12'habe, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9be, 12'hace, 12'hbde, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'hbbe, 12'haad, 12'h89b, 12'h67a, 12'h569, 12'h67a, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89c, 12'h88b, 12'h67a, 12'h469, 12'h67a, 12'h78b, 12'h78b, 12'h89c, 12'h9ac, 12'haad, 12'habd, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'habd, 12'hbcd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hbcd, 12'haac, 12'h9ac, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h88b, 12'h78a, 12'h77a, 12'h88a, 12'h99b, 12'habc, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'h9ac, 12'h99b, 12'haac, 12'habd, 12'haac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h779, 12'h678, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h777, 12'h777, 12'h777, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767, 12'h667, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h777, 12'h888, 12'h999, 12'hccc, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h777, 12'h444, 12'h444, 12'h444, 12'h344, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h334, 12'h334, 12'h335, 12'h345, 12'h345, 12'h456, 12'h457, 12'h568, 12'h579, 12'h67a, 12'h78a, 12'h78a, 12'h679, 12'h679, 12'h679, 12'h679, 12'h678, 12'h668, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h667, 12'h668, 12'h778, 12'h789, 12'h789, 12'h88a, 12'h89a, 12'h89a, 12'h899, 12'h889, 12'h789, 12'h678, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h678, 12'h778, 12'h778, 12'h778, 12'h789, 12'h88a, 12'h78a, 12'h78a, 12'h79b, 12'h89b, 12'h8ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 
12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h89d, 12'h89d, 12'h8ad, 12'h7ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 12'h7ad, 12'h48c, 12'h38c, 12'h7ae, 12'h8be, 12'h8bf, 12'h8be, 12'h8be, 12'h8be, 12'h7be, 12'h7ae, 12'h7ad, 12'h69d, 12'h58b, 12'h36a, 12'h459, 12'h359, 12'h359, 12'h56a, 12'h68b, 12'h79c, 12'h79c, 12'h8ac, 12'h9ad, 12'h9ac, 12'h67a, 12'h457, 12'h678, 12'haab, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddf, 12'habe, 12'h89d, 12'h89c, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hcce, 12'hace, 12'habe, 12'h9bd, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9be, 12'hace, 12'hbde, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 
12'hddd, 12'hddd, 12'hddd, 12'hcdd, 12'hccd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hbcc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hcdd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'hbce, 12'hbbe, 12'h9ac, 12'h89b, 12'h78b, 12'h67a, 12'h569, 12'h569, 12'h67a, 12'h78b, 12'h78a, 12'h67a, 12'h569, 12'h569, 12'h469, 12'h469, 12'h56a, 12'h78b, 12'h89c, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'haac, 12'habd, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbc, 12'haac, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h88b, 12'h88a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h99c, 12'h89b, 12'h89b, 12'h88b, 12'h78a, 12'h78a, 12'h88b, 12'h88b, 12'h99b, 12'haac, 12'hbbd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h789, 12'h778, 12'h667, 12'h556, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h767, 12'h667, 12'h666, 12'h666, 12'h666, 12'h667, 12'h777, 12'h778, 12'h888, 12'hbbb, 12'hdde, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h877, 12'h554, 12'h443, 12'h444, 12'h444, 12'h334, 12'h344, 12'h334, 12'h344, 12'h344, 12'h344, 12'h334, 12'h335, 12'h345, 12'h346, 12'h557, 12'h568, 12'h679, 12'h679, 12'h679, 12'h67a, 12'h679, 12'h679, 12'h568, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h678, 12'h778, 12'h789, 12'h88a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h889, 12'h789, 12'h678, 12'h567, 12'h667, 12'h657, 12'h657, 12'h667, 12'h667, 12'h678, 12'h668, 12'h778, 12'h779, 12'h789, 12'h78a, 12'h78a, 12'h78b, 12'h89b, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 
12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79d, 12'h89d, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 12'h9be, 12'h7ae, 12'h58d, 12'h49d, 12'h7ae, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8be, 12'h7be, 12'h7ae, 12'h7ad, 12'h69d, 12'h58c, 12'h36a, 12'h359, 12'h259, 12'h249, 12'h46a, 12'h78c, 12'h8ad, 12'h89c, 12'h89c, 12'h9ad, 12'h9ac, 12'h78a, 12'h358, 12'h778, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddf, 12'habe, 12'h89d, 12'h89c, 12'h9ad, 12'hbce, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9ad, 12'habd, 12'hbce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hddf, 12'hdef, 12'hddf, 12'hcdf, 12'hbce, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h79c, 12'h79c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9be, 12'hace, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 
12'hccc, 12'hccc, 12'hbbc, 12'hbbc, 12'hbbb, 12'hbbb, 12'hbbb, 12'habb, 12'haab, 12'haab, 12'haab, 12'haab, 12'haaa, 12'haaa, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'habb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbc, 12'hbbc, 12'hccc, 12'hccc, 12'hccc, 12'hcdd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccd, 12'hbcd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'hbbd, 12'hbce, 12'habd, 12'h9ac, 12'h89c, 12'h88b, 12'h67a, 12'h56a, 12'h569, 12'h569, 12'h569, 12'h569, 12'h569, 12'h569, 12'h67a, 12'h78b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ad, 
12'haad, 12'habd, 12'haad, 12'habd, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbbc, 12'haac, 12'h9ab, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h99b, 12'h88b, 12'h78a, 12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h88b, 12'h78b, 12'h88b, 12'h88b, 12'h78a, 12'h78a, 12'h89b, 12'h9ac, 12'habd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89a, 12'h778, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h766, 12'h766, 12'h777, 12'h777, 12'h777, 12'h888, 12'h99a, 12'hccd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'h888, 12'h555, 12'h443, 12'h444, 12'h444, 12'h344, 12'h344, 12'h334, 12'h334, 12'h344, 12'h345, 12'h335, 12'h335, 12'h346, 12'h457, 12'h568, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h668, 12'h568, 12'h568, 12'h568, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h678, 12'h678, 12'h778, 12'h789, 12'h88a, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h779, 12'h668, 12'h667, 12'h667, 12'h667, 12'h657, 12'h668, 12'h668, 12'h669, 12'h679, 12'h679, 12'h779, 12'h78a, 12'h78a, 12'h68a, 12'h79b, 12'h89b, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8bf, 12'h8bf, 12'h9be, 12'h9be, 12'h7ad, 12'h59c, 12'h69d, 12'h8be, 12'h9cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h69d, 12'h58c, 12'h47a, 12'h259, 12'h359, 12'h25a, 12'h47b, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9ac, 12'h68a, 12'h458, 12'h789, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdef, 12'hcdf, 12'habd, 12'habd, 12'habe, 12'habe, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'hbce, 12'hccf, 12'hcce, 12'hcdf, 12'hddf, 12'hdef, 12'hdef, 12'hddf, 12'hcde, 12'hbce, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ac, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9ce, 12'hbce, 12'hcde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hbbc, 12'hbbb, 
12'hbbb, 12'haab, 12'haab, 12'haaa, 12'haaa, 12'haaa, 12'h9aa, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'haaa, 12'haaa, 12'haaa, 12'haab, 12'haab, 12'habb, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hccd, 12'hccd, 12'hbbd, 12'habd, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'habd, 12'h9ac, 12'h99c, 12'h89b, 12'h78b, 12'h67a, 12'h569, 12'h67a, 12'h67a, 12'h67a, 12'h67a, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'hbcd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbbc, 12'h9ab, 12'h99b, 12'h89b, 12'h88a, 12'h78a, 12'h77a, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h89b, 12'h77a, 12'h78a, 12'h89b, 12'h99b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'haad, 12'habe, 12'hbbe, 12'habe, 12'habd, 12'haad, 12'h9ad, 12'h99c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h88b, 12'h88b, 12'h88b, 12'h78a, 12'h67a, 12'h67a, 12'h88b, 12'h9ac, 12'habd, 12'hbce, 
12'hcce, 12'hcce, 12'hcce, 12'hbce, 12'hbbe, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h88a, 12'h778, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h766, 12'h766, 12'h766, 12'h777, 12'h777, 12'h778, 12'h889, 12'hbbc, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddc, 12'h998, 12'h655, 12'h444, 12'h443, 12'h444, 12'h344, 12'h344, 12'h334, 12'h334, 12'h334, 12'h344, 12'h335, 12'h345, 12'h446, 12'h567, 12'h679, 12'h679, 12'h679, 12'h679, 12'h668, 12'h568, 12'h568, 12'h568, 12'h568, 12'h668, 12'h668, 12'h668, 12'h668, 12'h678, 12'h779, 12'h779, 12'h88a, 12'h89a, 12'h99b, 12'haab, 12'haab, 12'h9aa, 12'h99a, 12'h99a, 12'h99b, 12'h99b, 12'h99a, 12'h89a, 12'h89a, 12'h88a, 12'h789, 12'h678, 12'h668, 12'h658, 12'h668, 12'h668, 12'h779, 12'h77a, 12'h77a, 12'h67a, 12'h57a, 12'h67a, 12'h68a, 12'h68a, 12'h68b, 12'h78b, 12'h79b, 12'h79c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8bf, 12'h8bf, 12'h8bf, 12'h9cf, 12'h8be, 12'h7ad, 12'h59c, 12'h7ad, 12'h8be, 12'h9cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ad, 12'h69c, 12'h47b, 12'h25a, 12'h35a, 12'h46a, 12'h68c, 12'h8ad, 12'h9be, 12'h9ad, 12'h8ad, 12'h9bd, 12'h9ac, 12'h68a, 12'h458, 12'h889, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddf, 12'hcdf, 12'hcdf, 12'hace, 12'h9bd, 12'hbce, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'hcce, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hace, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h79c, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8bd, 12'h9bd, 12'hace, 12'hbde, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hccc, 12'hccc, 12'hbbc, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'haaa, 
12'h99a, 12'h999, 12'h999, 12'h899, 12'h889, 12'h889, 12'h889, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h889, 12'h889, 12'h889, 12'h889, 12'h889, 12'h889, 12'h889, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h99a, 12'h9aa, 12'haaa, 12'haab, 12'habb, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hccc, 12'hcdd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'hccd, 12'hbbd, 12'habd, 12'haac, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h89b, 12'h77a, 12'h77a, 12'h78b, 12'h89b, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habc, 12'hbcd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdee, 12'hccd, 12'hbbc, 12'haab, 12'h99b, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h89b, 12'h78a, 12'h779, 12'h789, 12'h88a, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'hbbe, 12'hbce, 12'hbbe, 12'habe, 12'haad, 12'h9ad, 12'h99c, 12'h89c, 12'h89c, 12'h89b, 12'h89c, 12'h99c, 12'h9ac, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h88b, 12'h78a, 12'h67a, 12'h67a, 12'h78a, 
12'h89b, 12'haac, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h78a, 12'h99c, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89a, 12'h789, 12'h778, 12'h777, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h567, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h766, 12'h776, 12'h777, 12'h777, 12'h788, 12'haaa, 12'hcdd, 12'hdee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h555, 12'h544, 12'h443, 12'h443, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h334, 12'h334, 12'h345, 12'h456, 12'h567, 12'h679, 12'h779, 12'h779, 12'h679, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h668, 12'h668, 12'h679, 12'h779, 12'h779, 12'h78a, 12'h89a, 12'h89a, 12'h9ab, 12'haab, 12'haab, 12'h9aa, 12'h99a, 12'h89a, 12'h99a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89a, 12'h89a, 12'h88a, 12'h779, 12'h668, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h89c, 12'h89d, 12'h89c, 12'h68b, 12'h57b, 12'h57b, 12'h58b, 12'h68b, 12'h68b, 12'h69b, 12'h79c, 12'h79c, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8bf, 12'h9bf, 12'h9cf, 12'h9ce, 12'h9be, 12'h7ad, 12'h69c, 12'h59d, 12'h7be, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7be, 12'h7ae, 12'h7ad, 12'h69d, 12'h48c, 12'h36b, 12'h36b, 12'h57b, 12'h79d, 12'h8ae, 12'h9be, 12'h9be, 12'h8ad, 12'h9bd, 12'h8ac, 12'h57a, 12'h568, 12'h99a, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdef, 12'hdef, 12'hdef, 12'hbcf, 12'habe, 12'hbce, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'habe, 12'hcdf, 12'hddf, 12'hddf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9ad, 12'h79c, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h9bd, 12'h9bd, 12'hbce, 12'hcde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbcc, 12'hbbc, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'haaa, 12'h99a, 12'h999, 12'h899, 12'h889, 
12'h888, 12'h788, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h778, 12'h677, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h788, 12'h788, 12'h888, 12'h889, 12'h889, 12'h889, 12'h899, 12'h999, 12'h99a, 12'h9aa, 12'haaa, 12'haab, 12'hbbb, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccd, 12'hbcd, 12'habd, 12'haac, 12'haad, 12'haac, 12'haad, 12'haad, 12'habd, 12'haad, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbce, 12'habd, 12'h99c, 12'h78b, 12'h89b, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hccd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccd, 12'habc, 12'h9ab, 12'h99b, 12'h89b, 12'h88a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h779, 12'h779, 12'h779, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'h9ad, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h89c, 12'h99c, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hbbd, 12'habd, 12'haad, 12'h89b, 12'h78b, 
12'h77a, 12'h67a, 12'h67a, 12'h78b, 12'h99b, 12'h9ac, 12'haac, 12'haad, 12'habd, 12'h99c, 12'h77a, 12'h88b, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h99c, 12'h99b, 12'h89b, 12'h89a, 12'h889, 12'h778, 12'h778, 12'h677, 12'h667, 12'h677, 12'h678, 12'h678, 12'h668, 12'h667, 12'h567, 12'h557, 12'h667, 12'h668, 12'h778, 12'h667, 12'h667, 12'h667, 12'h777, 12'h777, 12'h889, 12'hccc, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'haaa, 12'h655, 12'h544, 12'h443, 12'h443, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h334, 12'h334, 12'h345, 12'h456, 12'h567, 12'h678, 12'h779, 12'h679, 12'h668, 12'h568, 12'h558, 12'h558, 12'h568, 12'h668, 12'h779, 12'h779, 12'h789, 12'h78a, 12'h88a, 12'h89a, 12'h89a, 12'h99a, 12'h99a, 12'h9aa, 12'h99a, 12'h889, 12'h788, 12'h899, 12'h99a, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h88a, 12'h77a, 12'h669, 12'h569, 12'h67a, 12'h89c, 12'h9ad, 12'h9ae, 12'h9be, 12'h9be, 12'h8ad, 12'h69c, 12'h57b, 12'h47b, 12'h58b, 12'h68b, 12'h69c, 12'h79c, 12'h79c, 12'h89c, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ae, 12'h8be, 12'h8be, 12'h8ae, 12'h8bf, 12'h9bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9ce, 12'h8be, 12'h79d, 12'h69d, 12'h7ae, 12'h8be, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h7bf, 12'h7be, 12'h7be, 12'h7ae, 12'h7ae, 12'h69d, 12'h58c, 12'h47c, 12'h47c, 12'h68c, 12'h8ad, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9bd, 12'h89c, 12'h57a, 12'h569, 12'h9aa, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hdef, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'hbce, 12'hcdf, 12'hddf, 12'hcdf, 12'hbce, 12'hace, 12'habe, 12'habe, 12'habe, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h79c, 12'h79b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ac, 12'h9bd, 12'hacd, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbcc, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'haaa, 12'h99a, 12'h999, 12'h999, 12'h889, 12'h889, 12'h778, 12'h778, 12'h778, 
12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h566, 12'h566, 12'h566, 12'h567, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h677, 12'h778, 12'h778, 12'h778, 12'h788, 12'h888, 12'h889, 12'h889, 12'h999, 12'h99a, 12'h9aa, 12'haaa, 12'haab, 12'hbbb, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hcdd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hccd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 12'habd, 12'haad, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89c, 12'h99c, 12'h9ac, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'haad, 12'h9ad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'haad, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccd, 12'habc, 12'h9ab, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h779, 12'h779, 12'h789, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'h9ac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h99c, 12'h89c, 12'h88b, 12'h89b, 12'h89c, 12'h99c, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hcce, 12'hbce, 12'hbbe, 
12'habd, 12'h9ac, 12'h89b, 12'h77a, 12'h67a, 12'h77a, 12'h77a, 12'h88b, 12'h89b, 12'h78b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h789, 12'h778, 12'h778, 12'h677, 12'h678, 12'h778, 12'h779, 12'h779, 12'h779, 12'h679, 12'h679, 12'h78a, 12'h88a, 12'h89b, 12'h9ab, 12'h99b, 12'h89a, 12'h789, 12'h677, 12'h788, 12'hbbb, 12'hddd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'haaa, 12'h776, 12'h544, 12'h443, 12'h443, 12'h444, 12'h334, 12'h344, 12'h344, 12'h344, 12'h335, 12'h334, 12'h345, 12'h445, 12'h557, 12'h678, 12'h679, 12'h679, 12'h568, 12'h568, 12'h568, 12'h568, 12'h679, 12'h779, 12'h78a, 12'h78a, 12'h89a, 12'h89a, 12'h88a, 12'h88a, 12'h789, 12'h789, 12'h789, 12'h889, 12'h889, 12'h899, 12'h778, 12'h899, 12'haab, 12'habc, 12'habc, 12'haab, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h78a, 12'h679, 12'h56a, 12'h67b, 12'h89d, 12'h8ae, 12'h9bf, 12'h9cf, 12'h9cf, 12'h9bf, 12'h8ae, 12'h59c, 12'h48b, 12'h48b, 12'h68c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h89d, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ae, 12'h9ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8bf, 12'h9bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9be, 12'h8ae, 12'h79d, 12'h69d, 12'h79d, 12'h8be, 12'h9bf, 12'h8bf, 12'h8bf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h7bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h6ad, 12'h59d, 12'h48c, 12'h58c, 12'h69d, 12'h8ad, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h7ac, 12'h57a, 12'h679, 12'haab, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hdef, 12'hdef, 12'hcdf, 12'hcdf, 12'hddf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'hbce, 12'hcdf, 12'hbce, 12'hace, 12'habd, 12'h9bd, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79b, 12'h78a, 12'h78a, 12'h79b, 12'h89c, 12'h8ac, 12'h8ad, 12'h79b, 12'h78b, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9ac, 12'habc, 12'hccd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbcc, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'h9aa, 12'h99a, 12'h999, 12'h889, 12'h889, 12'h888, 12'h788, 12'h778, 12'h777, 12'h667, 12'h667, 12'h566, 
12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h567, 12'h667, 12'h667, 12'h667, 12'h677, 12'h778, 12'h778, 12'h778, 12'h788, 12'h788, 12'h889, 12'h889, 12'h999, 12'h99a, 12'h9aa, 12'haaa, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hcdd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'haad, 12'habe, 12'hbce, 12'hbce, 12'hbbe, 12'haad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccd, 12'habc, 12'haac, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h779, 12'h778, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h88a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h78b, 12'h88b, 12'h89b, 12'h89c, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 
12'hcce, 12'hbce, 12'hbbd, 12'haad, 12'h99c, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h789, 12'h678, 12'h677, 12'h667, 12'h678, 12'h789, 12'h88a, 12'h78a, 12'h78a, 12'h88a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'habd, 12'haac, 12'h88a, 12'h9aa, 12'hcdd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedd, 12'hbbb, 12'h877, 12'h554, 12'h443, 12'h443, 12'h443, 12'h334, 12'h334, 12'h344, 12'h344, 12'h345, 12'h334, 12'h345, 12'h445, 12'h556, 12'h567, 12'h668, 12'h668, 12'h568, 12'h568, 12'h568, 12'h679, 12'h78a, 12'h78a, 12'h89b, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h789, 12'h778, 12'h778, 12'h778, 12'h778, 12'h889, 12'h9aa, 12'h778, 12'h899, 12'hbbc, 12'hccd, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h88b, 12'h89b, 12'h78a, 12'h67a, 12'h57a, 12'h68c, 12'h8ae, 12'h8bf, 12'h9cf, 12'hacf, 12'hacf, 12'h9cf, 12'h9bf, 12'h7ad, 12'h58c, 12'h37b, 12'h68c, 12'h79d, 12'h79d, 12'h79d, 12'h79d, 12'h7ad, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8ae, 
12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8bf, 12'h8bf, 12'h9bf, 12'h9bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9be, 12'h7ae, 12'h79d, 12'h69d, 12'h79d, 12'h8ae, 12'h9bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h7ad, 12'h69d, 12'h58c, 12'h58c, 12'h69d, 12'h8ae, 12'h8be, 12'h8be, 12'h9be, 12'h9be, 12'h9ce, 12'h8ac, 12'h68a, 12'h78a, 12'hbbc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hdde, 12'hdef, 12'hdef, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'hbce, 12'hbcf, 12'habe, 12'h9ad, 12'h89c, 12'h78b, 12'h78a, 12'h9ac, 12'habd, 12'habd, 12'h9ad, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h79b, 12'h568, 12'h456, 12'h556, 12'h679, 12'h89c, 12'h8ac, 12'h8ac, 12'h78b, 12'h78b, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habc, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hbcc, 12'hbbb, 12'hbbb, 12'haab, 12'haaa, 12'h9aa, 12'h999, 12'h899, 12'h889, 12'h788, 12'h778, 12'h777, 12'h677, 12'h667, 12'h667, 12'h567, 12'h556, 12'h556, 12'h455, 12'h445, 
12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h566, 12'h566, 12'h667, 12'h667, 12'h667, 12'h677, 12'h777, 12'h778, 12'h778, 12'h788, 12'h888, 12'h889, 12'h999, 12'h99a, 12'h9aa, 12'haaa, 12'habb, 12'hbbb, 12'hbbb, 12'hccc, 12'hccc, 12'hcdd, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hcdd, 12'hbcd, 12'habc, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbce, 12'hbbe, 12'habd, 12'h9ad, 12'h89c, 12'h88c, 12'h99c, 12'haad, 12'habe, 12'habd, 12'h9ad, 12'h99c, 12'h89c, 12'h9ac, 12'haad, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habc, 12'hbcd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hccd, 12'haac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h778, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h768, 12'h778, 12'h778, 12'h769, 12'h669, 12'h779, 12'h88a, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h78b, 12'h78b, 12'h88b, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 
12'hcce, 12'hcce, 12'hcce, 12'hbbe, 12'habd, 12'h9ac, 12'h89b, 12'h88b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89a, 12'h889, 12'h778, 12'h678, 12'h668, 12'h668, 12'h779, 12'h88a, 12'h89a, 12'h89b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'haad, 12'habc, 12'hbbc, 12'hddd, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccb, 12'h988, 12'h555, 12'h544, 12'h443, 12'h443, 12'h333, 12'h334, 12'h334, 12'h344, 12'h345, 12'h335, 12'h345, 12'h445, 12'h446, 12'h457, 12'h567, 12'h568, 12'h568, 12'h669, 12'h679, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h78a, 12'h789, 12'h679, 12'h778, 12'h779, 12'h789, 12'h778, 12'h768, 12'h668, 12'h778, 12'h789, 12'h778, 12'h889, 12'hbbc, 12'hbbd, 12'hbbc, 12'haab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h67a, 12'h57b, 12'h69c, 12'h8ae, 12'h9cf, 12'h9cf, 12'h9cf, 12'hadf, 12'h9cf, 12'h9cf, 12'h8be, 12'h69d, 12'h38c, 12'h48c, 12'h69d, 12'h7ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 
12'h8bf, 12'h9bf, 12'h9bf, 12'h8bf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h8be, 12'h8be, 12'h8ae, 12'h79d, 12'h69d, 12'h79e, 12'h8ae, 12'h8bf, 12'h9bf, 12'h9bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h7ae, 12'h6ad, 12'h59d, 12'h59c, 12'h69d, 12'h8ae, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9bd, 12'h79b, 12'h89a, 12'hcdd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcde, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'habe, 12'hbce, 12'habd, 12'h89c, 12'h78a, 12'h557, 12'h445, 12'h567, 12'h89b, 12'habd, 12'h9ac, 12'h8ac, 12'h89c, 12'h89b, 12'h89c, 12'h89b, 12'h679, 12'h557, 12'h556, 12'h568, 12'h679, 12'h79c, 12'h89c, 12'h79c, 12'h78b, 12'h79b, 12'h79b, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hccd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbc, 12'hbbb, 12'haab, 12'haaa, 12'haaa, 12'h999, 12'h899, 12'h889, 12'h788, 12'h777, 12'h677, 12'h667, 12'h566, 12'h556, 12'h556, 12'h456, 12'h456, 12'h455, 12'h445, 12'h345, 12'h345, 12'h234, 
12'h234, 12'h234, 12'h234, 12'h134, 12'h134, 12'h234, 12'h234, 12'h335, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h567, 12'h667, 12'h667, 12'h667, 12'h677, 12'h778, 12'h778, 12'h788, 12'h888, 12'h889, 12'h899, 12'h99a, 12'h9aa, 12'haaa, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbbd, 12'haac, 12'h9ac, 12'haac, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'habd, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haad, 12'h89c, 12'h88c, 12'h88c, 12'h78b, 12'h78b, 12'h88c, 12'h89c, 12'h89c, 12'h88c, 12'h88c, 12'h88b, 12'h89c, 12'h9ad, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hbcd, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h778, 12'h778, 12'h678, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h779, 12'h779, 12'h678, 12'h679, 12'h779, 12'h88a, 12'h88a, 12'h78a, 12'h67a, 12'h77a, 12'h89b, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 
12'hbbe, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbd, 12'haad, 12'h99c, 12'h99c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h789, 12'h778, 12'h678, 12'h678, 12'h779, 12'h88a, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h99c, 12'hbbd, 12'hccd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'ha99, 12'h665, 12'h544, 12'h443, 12'h444, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h345, 12'h445, 12'h446, 12'h456, 12'h457, 12'h568, 12'h679, 12'h779, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h88a, 12'h78a, 12'h779, 12'h678, 12'h678, 12'h789, 12'h99a, 12'h88a, 12'h779, 12'h668, 12'h668, 12'h668, 12'h668, 12'h88a, 12'haac, 12'habc, 12'haac, 12'h9ac, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h78b, 12'h57a, 12'h47b, 12'h69c, 12'h7ae, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9df, 12'hacf, 12'h9cf, 12'h7be, 12'h59d, 12'h48c, 12'h48d, 12'h79e, 12'h8ae, 12'h9bf, 12'h8bf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9bf, 
12'h9bf, 12'h9cf, 12'h9cf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h8be, 12'h8be, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8bf, 12'h8bf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7bf, 12'h7ae, 12'h7ae, 12'h7ae, 12'h7ae, 12'h6ae, 12'h59d, 12'h69d, 12'h7ad, 12'h8be, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'hace, 12'h9bd, 12'h8ab, 12'habb, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hdde, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hcde, 12'hcde, 12'hbde, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'habd, 12'hbce, 12'h9bd, 12'h89c, 12'h78a, 12'h668, 12'h556, 12'h567, 12'h789, 12'h89b, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89c, 12'h78b, 12'h78a, 12'h679, 12'h679, 12'h67a, 12'h78b, 12'h79b, 12'h79b, 12'h78b, 12'h78b, 12'h79c, 12'h79c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hbcd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hbbc, 12'hbbb, 12'habb, 12'haaa, 12'h9aa, 12'h999, 12'h899, 12'h888, 12'h788, 12'h777, 12'h677, 12'h566, 12'h556, 12'h556, 12'h456, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h235, 12'h234, 12'h234, 
12'h234, 12'h124, 12'h124, 12'h124, 12'h124, 12'h134, 12'h234, 12'h234, 12'h344, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h667, 12'h667, 12'h677, 12'h778, 12'h788, 12'h788, 12'h889, 12'h899, 12'h999, 12'h99a, 12'haaa, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccd, 12'hbbd, 12'habc, 12'h9ac, 12'haac, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'habd, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h99c, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'haad, 12'h89c, 12'h78b, 12'h78b, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h77b, 12'h77b, 12'h77b, 12'h77b, 12'h88b, 12'h99c, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'hbcd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h779, 12'h779, 12'h778, 12'h679, 12'h679, 12'h679, 12'h679, 12'h669, 12'h78b, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 
12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'haad, 12'haac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h789, 12'h678, 12'h678, 12'h679, 12'h78a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h99b, 12'haac, 12'hbcd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbaa, 12'h777, 12'h555, 12'h444, 12'h444, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h445, 12'h446, 12'h446, 12'h457, 12'h568, 12'h679, 12'h78a, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h88a, 12'h78a, 12'h679, 12'h668, 12'h778, 12'h889, 12'haab, 12'haab, 12'h99a, 12'h779, 12'h668, 12'h668, 12'h679, 12'h89a, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h78b, 12'h57a, 12'h47b, 12'h69c, 12'h7ae, 12'h8bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8bf, 12'h6ae, 12'h59d, 12'h38c, 12'h58d, 12'h69d, 12'h8ae, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9cf, 
12'h9be, 12'h9be, 12'h9be, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8bf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h6ae, 12'h69d, 12'h59d, 12'h7ad, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'hace, 12'hace, 12'habd, 12'h9ab, 12'hbcc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hddf, 12'hdef, 12'hddf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hcce, 
12'hcce, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ad, 12'habd, 12'h9ad, 12'h89c, 12'h88b, 12'h78a, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h89b, 12'h79b, 12'h89b, 12'h79b, 12'h78b, 12'h79b, 12'h79b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hccc, 12'hbbb, 12'haab, 12'haaa, 12'h9aa, 12'h999, 12'h899, 12'h888, 12'h788, 12'h777, 12'h667, 12'h566, 12'h556, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h235, 12'h244, 12'h344, 12'h345, 12'h234, 12'h234, 12'h234, 12'h134, 
12'h124, 12'h024, 12'h024, 12'h024, 12'h024, 12'h134, 12'h134, 12'h234, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h456, 12'h556, 12'h556, 12'h566, 12'h667, 12'h677, 12'h677, 12'h778, 12'h778, 12'h788, 12'h888, 12'h889, 12'h999, 12'h99a, 12'haaa, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hccd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbcd, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'haac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h89c, 12'h78b, 12'h78b, 12'h78b, 12'h89c, 12'h9ac, 12'h9ad, 12'h9ac, 12'h88c, 12'h77b, 12'h67b, 12'h66b, 12'h77b, 12'h66b, 12'h77b, 12'h77b, 12'h77b, 12'h77b, 12'h77b, 12'h66b, 12'h77b, 12'h77b, 12'h77b, 12'h78b, 12'h89c, 12'haad, 12'haad, 12'haad, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h9ad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h88a, 12'h89a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h88a, 12'h779, 12'h779, 12'h778, 12'h778, 12'h779, 12'h779, 12'h779, 12'h778, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h679, 12'h679, 12'h679, 12'h78a, 12'h99c, 12'haad, 12'haad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 
12'hbbe, 12'hbbe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h789, 12'h678, 12'h678, 12'h789, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78b, 12'h88b, 12'h89b, 12'h99b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'haac, 12'hbcd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccb, 12'h988, 12'h665, 12'h444, 12'h444, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h445, 12'h446, 12'h446, 12'h457, 12'h568, 12'h679, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h78a, 12'h78a, 12'h779, 12'h679, 12'h779, 12'h88a, 12'h9ab, 12'haab, 12'h99b, 12'h88a, 12'h78a, 12'h67a, 12'h78a, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'h99c, 12'h9ac, 12'h89c, 12'h79c, 12'h78b, 12'h57a, 12'h47b, 12'h58c, 12'h7ad, 12'h8be, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h7bf, 12'h6ae, 12'h59d, 12'h48d, 12'h48d, 12'h59d, 12'h7ad, 12'h8ae, 12'h8be, 12'h8be, 12'h7ae, 
12'h7ad, 12'h7ae, 12'h7ae, 12'h7ae, 12'h8ae, 12'h8bf, 12'h9bf, 12'h9cf, 12'h9cf, 12'hacf, 12'hacf, 12'h9cf, 12'h9be, 12'h8be, 12'h8be, 12'h8bf, 12'h8cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h7ae, 12'h69d, 12'h59d, 12'h69d, 12'h8ad, 12'h9be, 12'h9be, 12'habe, 12'hace, 12'hacd, 12'habc, 12'hbbc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hcde, 12'hcdf, 12'hbcf, 12'hbce, 12'hace, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbde, 12'hbde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h78b, 12'h78b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hbce, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'h99a, 12'h999, 12'h899, 12'h888, 12'h778, 12'h677, 12'h667, 12'h566, 12'h456, 12'h445, 12'h345, 12'h344, 12'h334, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 
12'h134, 12'h134, 12'h134, 12'h134, 12'h134, 12'h134, 12'h234, 12'h244, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h445, 12'h445, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h667, 12'h667, 12'h677, 12'h777, 12'h778, 12'h778, 12'h788, 12'h888, 12'h889, 12'h999, 12'h9aa, 12'haaa, 12'habb, 12'hbbb, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h89b, 12'h78b, 12'h78b, 12'h67a, 12'h67a, 12'h78b, 12'h78b, 12'h77b, 12'h66a, 12'h56a, 12'h66a, 12'h66b, 12'h66a, 12'h55a, 12'h439, 12'h449, 12'h559, 12'h459, 12'h458, 12'h448, 12'h459, 12'h55a, 12'h66a, 12'h67b, 12'h78b, 12'h99c, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h99c, 12'h89c, 12'h89c, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'haad, 
12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'habc, 12'hbbd, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hbbc, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h88a, 12'h679, 12'h789, 12'h88a, 12'h89a, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h779, 12'h669, 12'h668, 12'h779, 12'h779, 12'h779, 12'h779, 12'h789, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h78a, 12'h88b, 12'h99c, 12'haad, 12'habd, 12'haad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 
12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h789, 12'h678, 12'h679, 12'h88a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h77a, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'haac, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'haaa, 12'h777, 12'h555, 12'h444, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h345, 12'h345, 12'h446, 12'h457, 12'h457, 12'h679, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h78a, 12'h78a, 12'h779, 12'h779, 12'h789, 12'h88a, 12'h89a, 12'h99b, 12'h99b, 12'h89b, 12'h78a, 12'h78a, 12'h78b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79b, 12'h57b, 12'h37a, 12'h58c, 12'h7ad, 12'h8be, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8bf, 12'h8bf, 12'h7ae, 12'h69e, 12'h48d, 12'h58d, 12'h69d, 12'h7ad, 12'h7ad, 12'h7ad, 12'h7ad, 
12'h7ae, 12'h7ae, 12'h8be, 12'h8bf, 12'h8bf, 12'h9cf, 12'h9cf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'h9cf, 12'h8be, 12'h8be, 12'h8bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h7ae, 12'h6ad, 12'h59d, 12'h69c, 12'h7ad, 12'h9be, 12'h9bd, 12'habd, 12'habd, 12'habc, 12'hbbc, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'hbcd, 12'hbcd, 12'habd, 12'habc, 12'h9ab, 12'habc, 12'hbce, 12'hbde, 12'hbde, 12'hbde, 12'hcde, 12'hcdf, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ac, 12'h99c, 12'h89c, 12'h9ac, 12'haad, 12'haad, 12'h9ad, 12'h89c, 12'h89c, 12'h89b, 12'h79b, 12'h79b, 12'h79c, 12'h79c, 12'h79b, 12'h79b, 12'h78b, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9cd, 12'hbde, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hbcc, 12'hbbb, 12'haab, 12'haaa, 12'h999, 12'h899, 12'h888, 12'h788, 12'h677, 12'h677, 12'h567, 12'h556, 12'h455, 12'h345, 12'h244, 12'h234, 12'h223, 12'h223, 12'h134, 12'h134, 12'h134, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 
12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h567, 12'h667, 12'h667, 12'h677, 12'h677, 12'h777, 12'h778, 12'h788, 12'h888, 12'h899, 12'h999, 12'haaa, 12'haab, 12'hbbb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h89c, 12'h9ac, 12'h9ad, 12'haad, 12'h9ac, 12'h89c, 12'h77b, 12'h67a, 12'h67b, 12'h77b, 12'h99d, 12'h99d, 12'h99d, 12'h98c, 12'h88c, 12'h66b, 12'h449, 12'h237, 12'h036, 12'h036, 12'h137, 12'h348, 12'h55a, 12'h56a, 12'h67a, 12'h78b, 12'h99c, 12'h9ac, 12'h89c, 12'h89b, 12'h78b, 12'h89b, 12'h89c, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'haad, 12'h9ad, 12'haad, 
12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'haad, 12'habd, 12'habc, 12'hbcd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdee, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h679, 12'h568, 12'h679, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h89b, 12'h88b, 12'h88a, 12'h88a, 12'h77a, 12'h77a, 12'h88a, 12'h88a, 12'h89b, 12'h99b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h89b, 12'h99c, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h789, 12'h779, 12'h78a, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78a, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'hbbd, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'h999, 12'h666, 12'h444, 12'h444, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h345, 12'h345, 12'h456, 12'h457, 12'h458, 12'h569, 12'h68a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h78a, 12'h78a, 12'h77a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h88b, 12'h88b, 12'h78b, 12'h78b, 12'h88b, 12'h79b, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h89c, 12'h79c, 12'h57b, 12'h37a, 12'h58c, 12'h6ad, 12'h8be, 12'h8bf, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h7ae, 12'h69e, 12'h69e, 12'h69e, 12'h7ae, 12'h8ae, 12'h8bf, 12'h8bf, 
12'h8bf, 12'h8bf, 12'h9cf, 12'h9cf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'h9cf, 12'h9bf, 12'h9be, 12'h9be, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7bf, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h6ad, 12'h59c, 12'h58c, 12'h69c, 12'h8ac, 12'h9bd, 12'h9bc, 12'habc, 12'habc, 12'hccd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hbbb, 12'haab, 12'hbce, 12'hbde, 12'hbde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hccf, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hbbc, 12'hbbb, 12'haaa, 12'h9aa, 12'h999, 12'h899, 12'h888, 12'h778, 12'h677, 12'h667, 12'h667, 12'h556, 12'h455, 12'h345, 12'h344, 12'h234, 12'h124, 12'h123, 12'h023, 12'h123, 12'h134, 12'h134, 12'h234, 12'h234, 12'h244, 12'h244, 12'h344, 12'h345, 12'h344, 12'h334, 
12'h234, 12'h234, 12'h244, 12'h244, 12'h244, 12'h244, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h345, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h567, 12'h667, 12'h667, 12'h667, 12'h677, 12'h677, 12'h777, 12'h778, 12'h788, 12'h889, 12'h999, 12'h9aa, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hccd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hccd, 12'hbbc, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'haad, 12'h99d, 12'h9ad, 12'haad, 12'hbbe, 12'hccf, 12'hcbf, 12'haae, 12'haae, 12'h99d, 12'h87c, 12'h77b, 12'h66b, 12'h77b, 12'h77b, 12'h77b, 12'h77b, 12'h66a, 12'h56a, 12'h66a, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h89c, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ad, 12'haad, 
12'haad, 12'h9ad, 12'h9ad, 12'h9ac, 12'haad, 12'habc, 12'habd, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdde, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h88a, 12'h568, 12'h457, 12'h668, 12'h779, 12'h779, 12'h78a, 12'h88a, 12'h88a, 12'h88b, 12'h88b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'haad, 
12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h779, 12'h789, 12'h89a, 12'h89b, 12'h89b, 12'h88a, 12'h77a, 12'h569, 12'h78b, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'hbcd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heed, 12'hccc, 12'h999, 12'h666, 12'h444, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h334, 12'h344, 12'h345, 12'h456, 12'h567, 12'h568, 12'h568, 12'h679, 12'h78a, 12'h88b, 12'h88b, 12'h89b, 12'h78b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h79c, 12'h67b, 12'h47a, 12'h58b, 12'h69d, 12'h8ae, 12'h8bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h7af, 12'h7ae, 12'h6ae, 12'h7ae, 12'h8bf, 12'h8bf, 12'h8bf, 
12'h9cf, 12'h9cf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'h9ce, 12'h9be, 12'h9be, 12'h9be, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7be, 12'h7ae, 12'h6ae, 12'h6ae, 12'h7ad, 12'h59c, 12'h48b, 12'h57a, 12'h79b, 12'h9ac, 12'habc, 12'hbbc, 12'hccd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haab, 12'habd, 12'hbdf, 12'hbde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hcce, 12'hccf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hace, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hbbc, 12'hbbb, 12'haaa, 12'h99a, 12'h899, 12'h889, 12'h788, 12'h777, 12'h677, 12'h667, 12'h566, 12'h456, 12'h455, 12'h345, 12'h244, 12'h234, 12'h134, 12'h123, 12'h123, 12'h123, 12'h023, 12'h134, 12'h134, 12'h134, 12'h234, 12'h244, 12'h344, 12'h345, 12'h344, 12'h244, 12'h244, 
12'h244, 12'h244, 12'h244, 12'h244, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h455, 12'h455, 12'h455, 12'h456, 12'h455, 12'h445, 12'h445, 12'h345, 12'h455, 12'h445, 12'h445, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h567, 12'h567, 12'h667, 12'h667, 12'h677, 12'h677, 12'h677, 12'h778, 12'h788, 12'h889, 12'h899, 12'h999, 12'haaa, 12'habb, 12'hbbb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbbc, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h99d, 12'h99d, 12'haae, 12'hbbe, 12'hbbf, 12'hbbe, 12'hbbe, 12'hbbe, 12'haae, 12'haae, 12'ha9e, 12'ha9d, 12'h99d, 12'haad, 12'haad, 12'h89c, 12'h78b, 12'h88b, 12'h99c, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ad, 
12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haac, 12'habd, 12'hbcd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdde, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h78a, 12'h457, 12'h346, 12'h668, 12'h779, 12'h779, 12'h779, 12'h78a, 12'h88a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h88b, 12'h88b, 12'h89b, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 
12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h789, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h679, 12'h669, 12'h77a, 12'h89b, 12'h9ad, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'haac, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h656, 12'h444, 12'h334, 12'h334, 12'h344, 12'h344, 12'h334, 12'h345, 12'h445, 12'h557, 12'h668, 12'h668, 12'h568, 12'h679, 12'h78a, 12'h88b, 12'h88b, 12'h89b, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h89b, 12'h89b, 12'h79b, 12'h79b, 12'h79b, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h67b, 12'h47b, 12'h58c, 12'h79d, 12'h7ae, 12'h8be, 12'h8bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h7af, 12'h6ae, 12'h6ae, 12'h7ae, 12'h7ae, 12'h8be, 
12'h9bf, 12'h9cf, 12'h9cf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hace, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7be, 12'h7ae, 12'h7ae, 12'h6ae, 12'h7ad, 12'h69c, 12'h47b, 12'h67a, 12'h9ab, 12'hbcc, 12'hddd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'habc, 12'hbce, 12'hbde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'hace, 12'hace, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hace, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hbbb, 12'habb, 12'haaa, 12'h999, 12'h899, 12'h888, 12'h778, 12'h677, 12'h667, 12'h566, 12'h556, 12'h455, 12'h345, 12'h345, 12'h234, 12'h134, 12'h134, 12'h034, 12'h134, 12'h134, 12'h134, 12'h034, 12'h034, 12'h134, 12'h234, 12'h244, 12'h244, 12'h344, 12'h345, 12'h344, 12'h344, 12'h344, 
12'h344, 12'h244, 12'h244, 12'h244, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h455, 12'h455, 12'h456, 12'h455, 12'h456, 12'h456, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h566, 12'h567, 12'h567, 12'h667, 12'h667, 12'h677, 12'h778, 12'h788, 12'h888, 12'h899, 12'h999, 12'h9aa, 12'haab, 12'hbbb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hbbc, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h99d, 12'h99d, 12'h99d, 12'ha9d, 12'haae, 12'haae, 12'haae, 12'hbae, 12'haae, 12'haae, 12'haae, 12'haae, 12'hbbe, 12'hcce, 12'haad, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h9ac, 12'haac, 12'habc, 12'habc, 12'hcde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdde, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h89a, 12'h568, 12'h447, 12'h789, 12'h889, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h77a, 12'h88b, 12'h88b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89b, 12'h88b, 12'h78b, 12'h88b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h77a, 12'h67a, 12'h67a, 12'h77a, 12'h88b, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h777, 12'h455, 12'h344, 12'h344, 12'h344, 12'h334, 12'h344, 12'h445, 12'h456, 12'h557, 12'h668, 12'h678, 12'h668, 12'h669, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h79b, 12'h79b, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h57a, 12'h47b, 12'h68c, 12'h79d, 12'h7ad, 12'h8ae, 12'h8bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8bf, 12'h7bf, 12'h7ae, 12'h6af, 12'h7ae, 12'h7ae, 12'h7ae, 
12'h8be, 12'h9bf, 12'h9cf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'hace, 12'hace, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7be, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ae, 12'h7ad, 12'h79c, 12'h68b, 12'h9ab, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'hbcd, 12'hbde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 12'hbce, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'hace, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hbce, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'haab, 12'h9aa, 12'h999, 12'h889, 12'h788, 12'h778, 12'h677, 12'h567, 12'h566, 12'h456, 12'h455, 12'h345, 12'h244, 12'h134, 12'h134, 12'h023, 12'h033, 12'h034, 12'h134, 12'h134, 12'h134, 12'h034, 12'h034, 12'h134, 12'h234, 12'h244, 12'h244, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 
12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h244, 12'h244, 12'h344, 12'h345, 12'h345, 12'h355, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h566, 12'h566, 12'h566, 12'h566, 12'h567, 12'h567, 12'h667, 12'h677, 12'h677, 12'h778, 12'h788, 12'h888, 12'h899, 12'h999, 12'h9aa, 12'haaa, 12'hbbb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hbbc, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99d, 12'h99d, 12'h99d, 12'h99d, 12'h99d, 12'haad, 12'haae, 12'haae, 12'haae, 12'ha9d, 12'ha9d, 12'ha9d, 12'h99d, 12'h99d, 12'h99c, 12'h89c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ad, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'hbcd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdde, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h9ac, 12'h88a, 12'h669, 12'h669, 12'h89a, 12'h99b, 12'haac, 12'h99b, 12'h88a, 12'h78a, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h77a, 12'h77a, 12'h88b, 12'h99c, 12'h9ac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78b, 12'h88b, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h89b, 12'h77a, 12'h77a, 12'h77a, 12'h78a, 12'h89b, 12'h9ac, 12'habd, 12'habe, 12'habd, 12'h9ac, 12'h99c, 12'h9ac, 12'hbbd, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'h999, 12'h666, 12'h445, 12'h444, 12'h444, 12'h344, 12'h445, 12'h455, 12'h556, 12'h556, 12'h668, 12'h778, 12'h679, 12'h669, 12'h679, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h89c, 12'h68b, 12'h57b, 12'h57b, 12'h68c, 12'h79d, 12'h79d, 12'h7ae, 12'h8bf, 12'h8bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9df, 12'h9df, 12'h9cf, 12'h9cf, 12'h8cf, 12'h7bf, 12'h7bf, 12'h7bf, 12'h8bf, 12'h8bf, 12'h7ae, 
12'h7ae, 12'h9be, 12'h9be, 12'h9ce, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7bf, 12'h7be, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ad, 12'h8ac, 12'h89b, 12'hbcc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'hbcd, 12'hbde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hbce, 12'hbce, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h9ad, 12'h9ad, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hbde, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hccd, 12'hccc, 12'hbbb, 12'haab, 12'h9aa, 12'h999, 12'h889, 12'h788, 12'h677, 12'h667, 12'h567, 12'h566, 12'h456, 12'h455, 12'h345, 12'h244, 12'h134, 12'h123, 12'h023, 12'h023, 12'h023, 12'h134, 12'h134, 12'h244, 12'h244, 12'h134, 12'h133, 12'h133, 12'h134, 12'h234, 12'h244, 12'h244, 12'h344, 12'h344, 12'h244, 12'h244, 
12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h244, 12'h244, 12'h244, 12'h244, 12'h344, 12'h345, 12'h345, 12'h355, 12'h455, 12'h455, 12'h456, 12'h566, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h566, 12'h567, 12'h567, 12'h667, 12'h667, 12'h677, 12'h677, 12'h778, 12'h788, 12'h788, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbc, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h99c, 12'h89c, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h99d, 12'h99d, 12'h99d, 12'h99d, 12'h99d, 12'h99d, 12'h99d, 12'h99d, 12'h88c, 12'h88c, 12'h88c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'hbcd, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdde, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h99b, 12'h88b, 12'h88a, 12'h88a, 12'h99b, 12'hbbc, 12'hbcd, 12'habc, 12'hbbc, 12'haac, 12'h89a, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h78a, 12'h88b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 
12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h88b, 12'h77a, 12'h77a, 12'h77a, 12'h88b, 12'h89c, 12'h9ac, 12'haad, 12'hbbe, 12'habd, 12'h99c, 12'h99c, 12'haad, 12'hcce, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h778, 12'h555, 12'h445, 12'h445, 12'h445, 12'h455, 12'h555, 12'h556, 12'h556, 12'h667, 12'h778, 12'h679, 12'h679, 12'h679, 12'h78a, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79b, 12'h78b, 12'h78b, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h89c, 12'h79b, 12'h68b, 12'h67b, 12'h68b, 12'h78c, 12'h79d, 12'h79d, 12'h7ae, 12'h8be, 12'h8bf, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9df, 12'h9df, 12'h9df, 12'h9cf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h9cf, 12'h8bf, 12'h8bf, 
12'h7ae, 12'h8be, 12'h9be, 12'h9be, 12'habe, 12'habe, 12'habe, 12'hace, 12'hace, 12'habe, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h7bf, 12'h7be, 12'h7be, 12'h7ae, 12'h7ae, 12'h7ad, 12'h8ac, 12'h9ac, 12'hcdd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbc, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'hace, 12'hace, 12'habe, 12'habe, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hcde, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hccd, 12'hccc, 12'hbbb, 12'haab, 12'h9aa, 12'h899, 12'h888, 12'h778, 12'h677, 12'h667, 12'h566, 12'h566, 12'h456, 12'h455, 12'h345, 12'h244, 12'h234, 12'h234, 12'h123, 12'h123, 12'h123, 12'h134, 12'h234, 12'h234, 12'h345, 12'h244, 12'h234, 12'h133, 12'h133, 12'h134, 12'h244, 12'h244, 12'h344, 12'h344, 12'h345, 12'h344, 12'h244, 
12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h244, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h455, 12'h455, 12'h456, 12'h556, 12'h566, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h677, 12'h677, 12'h678, 12'h778, 12'h778, 12'h788, 12'h789, 12'h889, 12'h99a, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hcdd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hddd, 12'hbbc, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h89c, 12'h99d, 12'h89c, 12'h88c, 12'h88c, 12'h88c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hbbc, 12'haab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'h9ac, 12'h99c, 12'h88b, 12'h88b, 12'h88b, 12'haac, 12'hccd, 12'hccd, 12'hccd, 12'hcde, 12'hbcd, 12'haab, 12'h88a, 12'h89a, 12'h89a, 12'h779, 12'h679, 12'h669, 12'h779, 12'h77a, 12'h88a, 12'h88b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h78b, 12'h88b, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 
12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h89c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h88b, 12'h89c, 12'h99c, 12'haad, 12'hbbe, 12'haad, 12'h99c, 12'haad, 12'hbbd, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'h999, 12'h666, 12'h444, 12'h445, 12'h445, 12'h455, 12'h455, 12'h556, 12'h556, 12'h567, 12'h778, 12'h779, 12'h679, 12'h569, 12'h67a, 12'h78b, 12'h89c, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h7ac, 12'h7ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ac, 12'h79c, 12'h68b, 12'h68b, 12'h68b, 12'h78c, 12'h79c, 12'h79c, 12'h69d, 12'h79d, 12'h7ae, 12'h8ae, 12'h8bf, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9df, 12'h9df, 12'h9df, 12'h9df, 12'h9df, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8bf, 
12'h8ae, 12'h8ae, 12'h9be, 12'h9be, 12'h9be, 12'habe, 12'habe, 12'habe, 12'habe, 12'habe, 12'hace, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h8ce, 12'h8ce, 12'h8bf, 12'h8bf, 12'h8be, 12'h8bf, 12'h8be, 12'h8bf, 12'h7be, 12'h7be, 12'h7ae, 12'h7ae, 12'h8ad, 12'h8ac, 12'h9ac, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbc, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'hace, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hace, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hcdd, 12'hccc, 12'hbbb, 12'haab, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h677, 12'h667, 12'h566, 12'h566, 12'h455, 12'h445, 12'h445, 12'h344, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h334, 12'h344, 12'h344, 12'h344, 12'h334, 12'h233, 12'h123, 12'h233, 12'h234, 12'h344, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h344, 
12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h345, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h456, 12'h456, 12'h566, 12'h566, 12'h567, 12'h556, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h889, 12'h99a, 12'h9aa, 12'habb, 12'hbbc, 12'hccc, 12'hcdd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'hddd, 12'habc, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78c, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'haac, 12'habc, 12'hccd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hbbc, 12'h9ab, 12'h9ab, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h88b, 12'h89b, 12'h99c, 12'habd, 12'hcce, 12'hdde, 12'hdde, 12'hccd, 12'habc, 12'h9ab, 12'hbbc, 12'hbbc, 12'h99b, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h779, 12'h77a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h78b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78b, 12'h77a, 12'h78b, 12'h88b, 12'h89c, 12'h9ac, 12'habd, 12'hbbe, 12'h9ad, 12'h9ac, 12'habd, 12'hcce, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h777, 12'h545, 12'h444, 12'h445, 12'h445, 12'h455, 12'h455, 12'h456, 12'h567, 12'h668, 12'h779, 12'h789, 12'h579, 12'h579, 12'h68a, 12'h89b, 12'h8ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79c, 12'h78b, 12'h68b, 12'h58b, 12'h68b, 12'h79c, 12'h8ac, 12'h79c, 12'h79c, 12'h69d, 12'h7ad, 12'h7ae, 12'h7be, 12'h7bf, 12'h8bf, 12'h8cf, 12'h9cf, 12'h9df, 12'h9df, 12'hadf, 12'hadf, 12'hadf, 12'h9cf, 12'h9cf, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9bf, 
12'h8be, 12'h8ae, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'habe, 12'hace, 12'hace, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h8ce, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h7be, 12'h7be, 12'h8be, 12'h8ae, 12'h8ad, 12'h8ac, 12'h9ac, 12'hcdd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbcc, 12'hbcd, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbcf, 12'hcce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'habe, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hbce, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haab, 12'haaa, 12'h999, 12'h889, 12'h788, 12'h777, 12'h667, 12'h666, 12'h566, 12'h555, 12'h455, 12'h445, 12'h445, 12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h334, 12'h223, 12'h123, 12'h233, 12'h334, 12'h344, 12'h445, 12'h455, 12'h445, 12'h445, 12'h445, 12'h344, 
12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h456, 12'h456, 12'h346, 12'h345, 12'h346, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h889, 12'h99a, 12'h9aa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbc, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h99c, 12'h89c, 12'h89b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h88b, 12'h89b, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'haac, 12'habc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hbbc, 12'h9ab, 12'h9ab, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h99c, 12'h88c, 12'h88b, 12'haad, 12'hcce, 12'hdde, 12'hcde, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'habc, 12'h89a, 12'h9ab, 12'haab, 12'h89a, 12'h779, 12'h779, 12'h779, 12'h779, 12'h78a, 12'h88a, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h99b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h89c, 12'h9ac, 12'haad, 12'hbbe, 12'habd, 12'h9ac, 12'haad, 12'hcce, 12'hdef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'h989, 12'h556, 12'h444, 12'h444, 12'h445, 12'h445, 12'h455, 12'h456, 12'h567, 12'h668, 12'h679, 12'h78a, 12'h579, 12'h579, 12'h57a, 12'h69b, 12'h79b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89b, 12'h79b, 12'h78b, 12'h78b, 12'h78b, 12'h79c, 12'h79c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h79c, 12'h79c, 12'h79d, 12'h7ad, 12'h8be, 12'h8be, 12'h8bf, 12'h8bf, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9df, 12'h9df, 12'hadf, 12'hadf, 12'h9cf, 12'h8cf, 12'h8cf, 12'h8cf, 12'h9cf, 12'h9bf, 12'h8be, 
12'h8be, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h8ce, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h7be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h89c, 12'h9ac, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbcc, 12'hbde, 12'hbde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habe, 12'hace, 12'hbce, 12'hbce, 12'hace, 12'habe, 12'habd, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h89c, 12'h88c, 12'h89c, 12'h89c, 12'h88b, 12'h79b, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ad, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hbcd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'habb, 12'haaa, 12'h999, 12'h889, 12'h788, 12'h677, 12'h667, 12'h566, 12'h556, 12'h556, 12'h455, 12'h455, 12'h445, 12'h445, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h444, 12'h444, 12'h344, 12'h344, 12'h344, 12'h344, 12'h334, 12'h233, 12'h123, 12'h233, 12'h344, 12'h344, 12'h445, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 
12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h456, 12'h456, 12'h566, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h346, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h467, 12'h467, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h789, 12'h889, 12'h99a, 12'h9aa, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'habc, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'haac, 12'habc, 12'hccd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hbcd, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89b, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'haad, 12'hbbd, 12'hcce, 12'hccd, 12'hcde, 12'hdee, 12'hdee, 12'hbcd, 12'habc, 12'hbcd, 12'hbcd, 12'h9ab, 12'h789, 12'h89a, 12'h89a, 12'h78a, 12'h779, 12'h679, 12'h779, 12'h88a, 12'h88a, 12'h88a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h67a, 12'h77a, 12'h78b, 12'h88b, 12'h89b, 12'h88b, 12'h88b, 12'h89c, 12'h99c, 12'haad, 12'hbbe, 12'hbbe, 12'h9ad, 12'h9ac, 12'hbbd, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'haaa, 12'h666, 12'h444, 12'h344, 12'h344, 12'h344, 12'h345, 12'h455, 12'h456, 12'h567, 12'h678, 12'h689, 12'h68a, 12'h57a, 12'h579, 12'h68a, 12'h79b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89b, 12'h79b, 12'h78b, 12'h78b, 12'h68b, 12'h68b, 12'h78b, 12'h79c, 12'h8ac, 12'h9ad, 12'h9bd, 12'h9bd, 12'h8ad, 12'h79c, 12'h79d, 12'h79d, 12'h7ae, 12'h8be, 12'h8be, 12'h8bf, 12'h8bf, 12'h8cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hadf, 12'hacf, 12'h9cf, 12'h9cf, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 
12'h8ad, 12'h8be, 12'h9be, 12'h9ce, 12'h9be, 12'h9be, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h8ac, 12'h9ac, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hddd, 12'hbbc, 12'hbce, 12'hbce, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 12'hbce, 12'hace, 12'habe, 12'habd, 12'habd, 12'hace, 12'hbce, 12'hace, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hace, 12'hbce, 12'hbce, 12'habe, 12'habd, 12'h9ad, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h88c, 12'h88b, 12'h88b, 12'h78b, 12'h88b, 12'h88b, 12'h78b, 12'h78b, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'habb, 12'h9aa, 12'h999, 12'h888, 12'h788, 12'h677, 12'h666, 12'h566, 12'h556, 12'h555, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h344, 12'h345, 12'h344, 12'h344, 12'h234, 12'h234, 12'h234, 12'h344, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 
12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h344, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h444, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h467, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h578, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h889, 12'h89a, 12'h9aa, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'haac, 12'h9ac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h99c, 12'h89c, 12'h89b, 12'h78b, 12'h78b, 12'h89b, 12'h88b, 12'h89b, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'habc, 12'hcdd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hddd, 12'hccd, 12'haab, 12'h99b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89c, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'ha9d, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'habd, 12'hbcd, 12'hcde, 12'hdee, 12'hcde, 12'hccd, 12'hcde, 12'hccd, 12'hbbc, 12'haac, 12'haab, 12'haac, 12'h99b, 12'h789, 12'h678, 12'h678, 12'h779, 12'h789, 12'h789, 12'h789, 12'h78a, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h669, 12'h569, 12'h669, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h89c, 12'haad, 12'hbbe, 12'hbbe, 12'haad, 12'h99c, 12'haad, 12'hcce, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h778, 12'h445, 12'h344, 12'h344, 12'h344, 12'h344, 12'h455, 12'h456, 12'h567, 12'h568, 12'h679, 12'h68a, 12'h78a, 12'h67a, 12'h57a, 12'h68a, 12'h78b, 12'h79b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h78b, 12'h78b, 12'h68b, 12'h68b, 12'h68b, 12'h78c, 12'h79c, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h7ad, 12'h79d, 12'h7ad, 12'h7ad, 12'h8be, 12'h8be, 12'h9bf, 12'h8bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hacf, 12'hacf, 12'hacf, 12'h9cf, 12'h9be, 12'h8be, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 
12'h8ad, 12'h8bd, 12'h9be, 12'h9ce, 12'h9ce, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h8ad, 12'habd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbcc, 12'hbcd, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcdf, 12'hcdf, 12'hcdf, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcdf, 12'hcce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habe, 12'habe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habe, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h89c, 12'h88c, 12'h88b, 12'h88b, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h79b, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hace, 12'hbcd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haab, 12'h9aa, 12'h899, 12'h888, 12'h777, 12'h677, 12'h666, 12'h556, 12'h555, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h344, 12'h334, 12'h334, 12'h344, 12'h345, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 
12'h345, 12'h344, 12'h344, 12'h345, 12'h445, 12'h445, 12'h445, 12'h344, 12'h234, 12'h234, 12'h334, 12'h344, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h889, 12'h89a, 12'h9aa, 12'hbbb, 12'hbbc, 12'hccc, 12'hcdd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 
12'hbcd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hddd, 12'hccd, 12'haab, 12'h99b, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'ha9d, 12'ha9d, 12'ha9d, 12'h99d, 12'h99c, 12'h89c, 12'h9ac, 12'habd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hbcd, 12'hbbd, 12'habc, 12'haac, 12'h99b, 12'h88a, 12'h889, 12'h889, 12'h789, 12'h779, 12'h668, 12'h678, 12'h679, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h78a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h679, 12'h458, 12'h679, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h89c, 12'h9ac, 12'haad, 12'hbbe, 12'habe, 12'h9ad, 12'h99c, 12'h9ac, 12'hbbe, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h999, 12'h556, 12'h344, 12'h444, 12'h344, 12'h344, 12'h345, 12'h456, 12'h567, 12'h567, 12'h568, 12'h779, 12'h78a, 12'h78a, 12'h67a, 12'h67a, 12'h68a, 12'h68a, 12'h68b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h68b, 12'h68b, 12'h68b, 12'h78b, 12'h79c, 12'h89c, 12'h89d, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 12'h7ad, 12'h8ae, 12'h8be, 12'h9bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hacf, 12'hacf, 12'hacf, 12'hacf, 12'h9ce, 12'h9bd, 12'h8ad, 12'h7ac, 12'h7ac, 12'h79c, 12'h79c, 
12'h7ad, 12'h8bd, 12'h9be, 12'h9be, 12'h9be, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h8ad, 12'hbbd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbc, 12'hbce, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hcdf, 12'hcdf, 12'hcdf, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'h9ad, 12'h89c, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78a, 12'h78b, 12'h78b, 12'h89b, 12'h8ac, 12'h7ac, 12'h79c, 12'h79b, 12'h7ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hace, 12'hbcd, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'habb, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h667, 12'h666, 12'h556, 12'h455, 12'h455, 12'h445, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h344, 12'h234, 12'h234, 12'h234, 12'h344, 12'h345, 12'h345, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h668, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h889, 12'h99a, 12'haab, 12'hbbb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'hbcd, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hddd, 12'hccd, 12'haac, 12'h99b, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'ha9d, 12'ha9d, 12'haad, 12'h9ad, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'haac, 12'hbbd, 12'hbcd, 12'haac, 12'habc, 12'habc, 12'haac, 12'h89b, 12'h78a, 12'h88a, 12'h89a, 12'h889, 12'h668, 12'h568, 12'h568, 12'h457, 12'h458, 12'h78a, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h88b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h78a, 12'h89b, 12'h9ac, 12'h99c, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habe, 12'haad, 12'h99c, 12'h89c, 12'h9ac, 12'hbbd, 12'hcce, 12'hdde, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h778, 12'h445, 12'h444, 12'h344, 12'h344, 12'h345, 12'h456, 12'h567, 12'h567, 12'h568, 12'h679, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h68a, 12'h68a, 12'h78b, 12'h68b, 12'h68b, 12'h68b, 12'h68b, 12'h78c, 12'h79c, 12'h79c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 12'h8ae, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9cf, 12'hacf, 12'hacf, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h8ad, 12'h7ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 
12'h7ad, 12'h8bd, 12'h8bd, 12'h8be, 12'h9bd, 12'h8bd, 12'h9bd, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h9bd, 12'hbcd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hccd, 12'hbce, 12'hbde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 
12'hbde, 12'hcde, 12'hcde, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'habd, 12'h9ac, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h77a, 12'h77a, 12'h77a, 12'h77b, 12'h77b, 12'h87b, 12'h78b, 12'h77b, 12'h77b, 12'h77b, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h78a, 12'h78a, 12'h77a, 12'h78a, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hcdd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h667, 12'h566, 12'h556, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 12'h345, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h445, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h344, 12'h234, 12'h234, 12'h234, 12'h344, 12'h345, 12'h345, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h566, 12'h567, 12'h567, 12'h466, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h889, 12'h99a, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'habd, 12'hbbe, 12'hbbd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'hbbd, 12'hdde, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hdde, 12'hccd, 12'habc, 12'h99b, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88b, 12'h88b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99d, 12'haad, 12'haad, 12'haad, 12'haad, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h88b, 12'h78a, 12'h88a, 12'h88a, 12'h779, 12'h668, 12'h678, 12'h678, 12'h568, 12'h458, 12'h77a, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 
12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h99b, 12'h99c, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'h9ac, 12'h89c, 12'h99c, 12'haad, 12'hbbd, 12'hbcd, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'h9aa, 12'h666, 12'h445, 12'h344, 12'h344, 12'h345, 12'h455, 12'h456, 12'h557, 12'h557, 12'h568, 12'h679, 12'h78a, 12'h78b, 12'h78b, 12'h89b, 12'h89b, 12'h79b, 12'h79c, 12'h79c, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 12'h8ad, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'hace, 12'hace, 12'hace, 12'hace, 12'hace, 12'h9bd, 12'h9ad, 12'h8ac, 12'h89c, 12'h79c, 12'h79c, 12'h7ac, 12'h7ac, 
12'h8ad, 12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ad, 12'h9bd, 12'hcce, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hcdd, 12'hbce, 12'hbce, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 
12'hbde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bc, 12'h9bd, 12'habd, 12'hbce, 12'habd, 12'h89c, 12'h78b, 12'h78a, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h67a, 12'h67a, 12'h67a, 12'h67a, 12'h679, 12'h679, 12'h67a, 12'h67a, 12'h68a, 12'h79b, 12'h79b, 12'h7ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hbcd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h667, 12'h566, 12'h556, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h445, 
12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h344, 12'h134, 12'h234, 12'h234, 12'h334, 12'h344, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h899, 12'h99a, 12'haab, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hcde, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'hccd, 12'heef, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hdde, 12'hccd, 12'hbbc, 12'h9ab, 12'h99b, 12'h99b, 12'h99c, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'haad, 12'haad, 12'haad, 12'haad, 12'h9ad, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h89b, 12'h88b, 12'h88a, 12'h88a, 12'h89b, 12'h89b, 12'h9ab, 12'h89b, 12'h88b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h89b, 12'h99c, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccc, 12'h889, 12'h566, 12'h445, 12'h344, 12'h344, 12'h445, 12'h456, 12'h456, 12'h457, 12'h458, 12'h569, 12'h57a, 12'h78a, 12'h79b, 12'h89b, 12'h79c, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h7ac, 12'h7ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9be, 12'habe, 12'habe, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ac, 12'h89c, 12'h89c, 12'h7ac, 12'h79c, 12'h7ac, 12'h8ad, 
12'h8ad, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8bd, 12'h8ad, 12'habd, 12'hcde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hcce, 12'hbce, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 
12'hbde, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hacd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h77b, 12'h77b, 12'h77b, 12'h78b, 12'h88b, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h88b, 12'h78b, 12'h77a, 12'h77a, 12'h67a, 12'h78a, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h79c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'hacd, 12'hbcd, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'hddd, 12'hccd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h667, 12'h566, 12'h456, 12'h455, 12'h455, 12'h445, 12'h345, 12'h445, 12'h445, 12'h455, 12'h455, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h445, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h234, 12'h234, 12'h234, 12'h234, 12'h244, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h889, 12'h899, 12'h99a, 12'haab, 12'habb, 12'hbbc, 12'hccc, 12'hcdd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'heff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'h9ac, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'haad, 12'habd, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbe, 12'habe, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'habc, 12'hdde, 12'heef, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hddd, 12'hccd, 12'hbbc, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h88a, 12'h78a, 12'h88a, 12'h88a, 12'h88b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h89c, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habd, 12'h9ac, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h78a, 12'h88b, 12'h89b, 12'h89c, 12'h99c, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'habd, 12'hbbd, 12'habc, 12'habc, 12'hbbc, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'h888, 12'h666, 12'h455, 12'h444, 12'h345, 12'h345, 12'h446, 12'h457, 12'h458, 12'h569, 12'h569, 12'h67a, 12'h78b, 12'h79b, 12'h79c, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ac, 12'h79c, 12'h79c, 12'h79c, 12'h8ac, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 
12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8bd, 12'h9bd, 12'habd, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbcd, 12'hbce, 12'hcce, 12'hcde, 12'hbde, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h88b, 12'h99c, 12'h99c, 12'haad, 12'haad, 12'haad, 12'h99d, 12'h99c, 12'h99c, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h88c, 12'h89c, 12'h99c, 12'h99c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'hbcd, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haab, 12'h999, 12'h889, 12'h778, 12'h677, 12'h566, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h566, 12'h556, 12'h556, 12'h456, 12'h455, 12'h355, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h445, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h244, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h455, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h789, 12'h889, 12'h89a, 12'h99a, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbbd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'hccd, 12'heef, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hddd, 12'hcdd, 12'hbbc, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h99b, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h89a, 12'h78a, 12'h78a, 12'h88a, 12'h78a, 12'h88a, 12'h88b, 12'h98b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h88c, 12'h88b, 12'h89b, 12'h89c, 12'h89c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habd, 12'habc, 12'h9ab, 12'h9ab, 12'hbbc, 12'hbcc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'haab, 12'h888, 12'h666, 12'h455, 12'h445, 12'h445, 12'h446, 12'h456, 12'h568, 12'h569, 12'h67a, 12'h68b, 12'h78b, 12'h79b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ac, 12'h7ac, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 
12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8bd, 12'h9bd, 12'hacd, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bc, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h79b, 12'h78a, 12'h89b, 12'h88b, 12'h89b, 12'h99c, 12'haac, 12'haad, 12'hbbd, 12'hbad, 12'haad, 12'haad, 12'haad, 12'h99d, 12'h99c, 12'h99c, 12'h99c, 12'h88c, 12'h88c, 12'h88c, 12'h89c, 12'h89c, 12'h88c, 12'h88c, 12'h88c, 12'h88b, 12'h88b, 12'h78b, 12'h88b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9bc, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'hacd, 12'hbde, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hccc, 12'hbbc, 12'haab, 12'h99a, 12'h889, 12'h788, 12'h677, 12'h567, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h345, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h244, 12'h234, 12'h234, 12'h234, 12'h134, 12'h234, 12'h245, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h345, 12'h345, 12'h345, 12'h235, 12'h345, 12'h445, 12'h455, 12'h445, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h789, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hdde, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habc, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hcdd, 12'hbbc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h88a, 12'h88a, 12'h789, 12'h789, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'h9ad, 12'haad, 12'h9ad, 12'haad, 12'habd, 12'habc, 12'haab, 12'h89a, 12'h889, 12'h9aa, 12'hbbc, 12'hccc, 12'hddd, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccd, 12'haaa, 12'h888, 12'h666, 12'h555, 12'h445, 12'h346, 12'h357, 12'h569, 12'h78a, 12'h79b, 12'h79b, 12'h79b, 12'h79b, 12'h79c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8be, 
12'h9be, 12'h9bf, 12'h9bf, 12'h9be, 12'h9be, 12'h8be, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h79c, 12'h79c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'habd, 12'hbce, 12'hcde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hcdd, 12'hbcd, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bc, 12'h9ac, 12'h8ab, 12'h89b, 12'h8ab, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'haad, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h98c, 12'h99c, 12'h88c, 12'h88c, 12'h88c, 12'h88b, 12'h88b, 12'h88c, 12'h88c, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'hbce, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hccc, 12'hbbc, 12'haab, 12'h99a, 12'h899, 12'h788, 12'h677, 12'h567, 12'h556, 12'h456, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h566, 12'h556, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h245, 12'h234, 12'h244, 12'h244, 12'h245, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h445, 12'h345, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h234, 12'h234, 12'h134, 12'h134, 12'h234, 12'h235, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h245, 12'h345, 12'h445, 12'h455, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h355, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h457, 12'h457, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h568, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h789, 12'h789, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbcd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'hcde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hddd, 12'hcdd, 12'hbbc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h88a, 12'h88a, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h88b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'haac, 12'h99b, 12'h789, 12'h788, 12'h999, 12'habb, 12'hbcc, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h667, 12'h456, 12'h456, 12'h356, 12'h568, 12'h78a, 12'h89b, 12'h89c, 12'h79c, 12'h79b, 12'h79c, 12'h79c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8be, 12'h9be, 
12'h9be, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9ce, 12'h9be, 12'h8ad, 12'h8ac, 12'h79c, 12'h79b, 12'h68b, 12'h69b, 12'h79c, 12'h7ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'hbce, 12'hddf, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbcd, 12'hbce, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hace, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h78b, 12'h77b, 12'h77b, 12'h77b, 12'h78b, 12'h78b, 12'h78b, 12'h78a, 12'h78a, 12'h78b, 12'h78b, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bd, 12'habd, 12'habd, 12'hbcd, 12'hcde, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hccc, 12'hbcc, 12'habb, 12'h9aa, 12'h899, 12'h888, 12'h778, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h556, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h245, 12'h235, 12'h234, 12'h234, 12'h234, 12'h235, 12'h245, 12'h345, 12'h345, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h235, 12'h234, 12'h134, 12'h134, 12'h134, 12'h235, 12'h245, 12'h345, 12'h456, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h245, 12'h345, 12'h445, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h457, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h667, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h788, 12'h789, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'habb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 
12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbbe, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'hccd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hcdd, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h89b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'h9ab, 12'h88a, 12'h789, 12'h788, 12'h889, 12'h9aa, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'haaa, 12'h888, 12'h667, 12'h556, 12'h457, 12'h458, 12'h679, 12'h89b, 12'h8ac, 12'h89c, 12'h79b, 12'h79b, 12'h79c, 12'h89c, 12'h79c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h89c, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9be, 12'h9be, 
12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8bd, 12'h8ad, 12'h89c, 12'h79c, 12'h78c, 12'h68b, 12'h58b, 12'h68b, 12'h69c, 12'h7ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9bd, 12'h9be, 12'h9be, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'hace, 12'hcde, 12'hdef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hbcd, 12'hbcd, 12'hbce, 
12'hbce, 12'hbce, 12'hbce, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78b, 12'h78b, 12'h88b, 12'h78b, 12'h78b, 12'h78b, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hcde, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbcc, 12'hbbb, 12'haaa, 12'h999, 12'h889, 12'h778, 12'h667, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h245, 12'h234, 12'h234, 12'h235, 12'h234, 12'h234, 12'h235, 12'h345, 12'h345, 12'h346, 12'h345, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h346, 12'h345, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h234, 12'h134, 12'h134, 12'h134, 12'h235, 12'h245, 12'h345, 12'h346, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h778, 12'h788, 12'h789, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'hbbb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 
12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'hbbd, 12'hcdd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hcdd, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h78a, 12'h88a, 12'h88a, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h889, 12'h899, 12'haab, 12'hbcc, 12'hccc, 12'hddd, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccc, 12'habb, 12'h889, 12'h777, 12'h557, 12'h567, 12'h679, 12'h89b, 12'h8ac, 12'h8ac, 12'h79c, 12'h79b, 12'h79b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h79c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 
12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h79d, 12'h79c, 12'h68c, 12'h68c, 12'h68b, 12'h68c, 12'h69c, 12'h79c, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9be, 12'h9be, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'habd, 12'hbce, 12'hcde, 12'hdef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbcd, 12'hbcd, 12'hbcd, 
12'hbce, 12'hbce, 12'hbce, 12'hacd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bd, 12'h9ac, 12'h8ac, 12'h89c, 12'h89b, 12'h89b, 12'h78b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78b, 12'h79b, 12'h79b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bd, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hcdd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hccd, 12'hbcc, 12'hbbb, 12'haaa, 12'h99a, 12'h889, 12'h788, 12'h677, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h245, 12'h235, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h235, 12'h345, 12'h345, 12'h346, 12'h346, 12'h356, 12'h456, 12'h456, 12'h456, 12'h356, 12'h346, 12'h346, 
12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h346, 12'h345, 12'h345, 12'h245, 12'h235, 12'h235, 12'h134, 12'h134, 12'h235, 12'h245, 12'h345, 12'h345, 12'h346, 12'h456, 12'h446, 12'h346, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h778, 12'h788, 12'h788, 12'h889, 12'h889, 12'h999, 12'h9aa, 12'haab, 12'hbbb, 12'hbcc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 
12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hccd, 12'h9ac, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'hbbd, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hcdd, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h78a, 12'h78a, 12'h79a, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h889, 12'h889, 12'h899, 12'h9aa, 12'hbbb, 12'hccc, 12'hcdd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccd, 12'hbbb, 12'h889, 12'h678, 12'h567, 12'h679, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79c, 12'h79b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 
12'h7ad, 12'h79d, 12'h79d, 12'h79d, 12'h79d, 12'h79c, 12'h78c, 12'h78c, 12'h68c, 12'h68c, 12'h68c, 12'h79c, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 12'hbce, 12'hcde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hccd, 12'hbcd, 12'hbcd, 
12'hbcd, 12'hbcd, 12'hbcd, 12'hacd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78b, 12'h78b, 12'h88b, 12'h89b, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'hacd, 12'hacd, 12'hbcd, 12'hbcd, 12'hcde, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hccd, 12'hbcc, 12'habb, 12'haaa, 12'h99a, 12'h889, 12'h788, 12'h677, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h566, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h235, 12'h234, 12'h234, 12'h234, 12'h235, 12'h345, 12'h345, 12'h346, 12'h346, 12'h456, 12'h456, 12'h456, 12'h456, 12'h356, 12'h456, 12'h446, 
12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h345, 12'h345, 12'h245, 12'h235, 12'h235, 12'h235, 12'h235, 12'h235, 12'h245, 12'h345, 12'h345, 12'h345, 12'h346, 12'h446, 12'h446, 12'h346, 12'h346, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h467, 12'h457, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h788, 12'h789, 12'h889, 12'h889, 12'h899, 12'h9aa, 12'haaa, 12'hbbb, 12'hccc, 12'hcdd, 12'hddd, 12'hdee, 12'heee, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdee, 12'hbbd, 12'h9ac, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habc, 12'hccd, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hddd, 12'hbcc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h899, 12'h99a, 12'haab, 12'hbcc, 12'hccd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h889, 12'h678, 12'h679, 12'h89a, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h79b, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h79c, 12'h79c, 
12'h79d, 12'h79d, 12'h89d, 12'h89d, 12'h89d, 12'h89d, 12'h89d, 12'h79d, 12'h79d, 12'h78d, 12'h79d, 12'h8ad, 12'h8ad, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 12'hbce, 12'hddf, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hcdd, 12'hcde, 12'hbcd, 
12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h79b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcde, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbcc, 12'hbbb, 12'haaa, 12'h99a, 12'h889, 12'h788, 12'h678, 12'h667, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h556, 12'h456, 12'h456, 12'h355, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h235, 12'h234, 12'h234, 12'h234, 12'h345, 12'h345, 12'h346, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h346, 12'h346, 12'h346, 12'h346, 12'h456, 12'h456, 12'h456, 12'h346, 12'h345, 12'h345, 12'h245, 12'h245, 12'h235, 12'h235, 12'h235, 12'h235, 12'h245, 12'h245, 12'h345, 12'h345, 12'h346, 12'h346, 12'h456, 12'h456, 12'h456, 12'h346, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h455, 12'h455, 12'h456, 12'h455, 12'h456, 12'h456, 12'h456, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h668, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h788, 12'h788, 12'h789, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbcd, 12'h9ab, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h9ac, 12'h9ac, 12'haac, 12'haad, 12'habd, 12'haad, 12'haac, 12'haac, 12'haad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'hdde, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hddd, 12'hbcc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89b, 12'h88a, 12'h88a, 12'h88a, 12'h78a, 12'h78a, 12'h88a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h99b, 12'h99b, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'haaa, 12'hbbb, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'habb, 12'h889, 12'h789, 12'h88a, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h79b, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h89c, 12'h89c, 12'h79c, 12'h78c, 12'h78d, 
12'h79d, 12'h89d, 12'h89e, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h79d, 12'h79d, 12'h79d, 12'h7ad, 12'h8bd, 12'h8be, 12'h9be, 12'h9be, 12'h8be, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'habd, 12'hcde, 12'hdef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hcde, 12'hcde, 
12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'habd, 12'habd, 12'habc, 12'h9bc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'hbcd, 12'hbcd, 12'hccd, 12'hcde, 12'hcde, 12'hdee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbc, 12'hbbb, 12'haaa, 12'h99a, 12'h889, 12'h788, 12'h678, 12'h667, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h234, 12'h234, 12'h234, 12'h345, 12'h346, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h346, 12'h446, 12'h346, 12'h446, 12'h456, 12'h456, 12'h456, 12'h346, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h235, 12'h235, 12'h235, 12'h245, 12'h245, 12'h345, 12'h345, 12'h345, 12'h346, 12'h356, 12'h456, 12'h456, 12'h456, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h678, 12'h778, 12'h778, 12'h778, 12'h788, 12'h789, 12'h889, 12'h999, 12'h9aa, 12'habb, 12'hbcc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'hccd, 12'haac, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'haac, 12'hbcd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hddd, 12'hbcd, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'haab, 12'haab, 12'haaa, 12'haab, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hcdd, 12'habb, 12'h89a, 12'h89a, 12'h89a, 12'h9ab, 12'h9ac, 12'habc, 12'h9ac, 12'h89b, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h78c, 12'h78c, 12'h78c, 12'h78d, 
12'h89e, 12'h9ae, 12'h9af, 12'h9bf, 12'h9bf, 12'h9af, 12'h9ae, 12'h8ae, 12'h7ae, 12'h79d, 12'h7ad, 12'h7ad, 12'h8be, 12'h8be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8bd, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h9ad, 12'h9bd, 12'hbce, 12'hcde, 12'hdef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hdee, 12'hcde, 
12'hcce, 12'hbcd, 12'hbcd, 12'hacd, 12'habd, 12'habd, 12'habc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'hbcd, 12'hccd, 12'hcde, 12'hdde, 12'hdee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haab, 12'haaa, 12'h99a, 12'h889, 12'h788, 12'h678, 12'h667, 12'h567, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h235, 12'h234, 12'h234, 12'h235, 12'h345, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h346, 12'h346, 12'h346, 12'h346, 12'h456, 12'h456, 12'h346, 12'h346, 12'h345, 12'h345, 12'h245, 12'h235, 12'h235, 12'h235, 12'h245, 12'h245, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h346, 12'h456, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h677, 12'h677, 12'h677, 12'h677, 12'h678, 12'h678, 12'h778, 12'h788, 12'h889, 12'h899, 12'h99a, 12'haaa, 12'hbbb, 12'hccc, 12'hccd, 12'hddd, 12'hdde, 
12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hbbc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'habc, 12'hbcd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hbcd, 12'habc, 12'haac, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'haab, 12'haab, 12'habb, 12'hbbb, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hccd, 12'habb, 12'h99a, 12'h89a, 12'h89b, 12'h9ab, 12'h9ac, 12'h9ac, 12'h89b, 12'h79b, 12'h79b, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 12'h78c, 12'h78c, 12'h78c, 12'h78c, 12'h78c, 12'h78d, 12'h88d, 12'h89e, 
12'h9ae, 12'h9bf, 12'h9bf, 12'habf, 12'h9bf, 12'h9af, 12'h8ae, 12'h8ae, 12'h8ae, 12'h7ad, 12'h7ad, 12'h7ad, 12'h8be, 12'h8be, 12'h8be, 12'h9be, 12'h8be, 12'h8be, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'habd, 12'hbce, 12'hcde, 12'hdef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdef, 12'hdde, 
12'hcde, 12'hcce, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9ac, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h78b, 12'h89b, 12'h89b, 12'h8ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89b, 12'h89c, 12'h89b, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hdde, 12'hdee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hccd, 12'hccc, 12'hbbb, 12'haab, 12'h99a, 12'h999, 12'h889, 12'h778, 12'h677, 12'h667, 12'h566, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h235, 12'h235, 12'h235, 12'h235, 12'h245, 12'h345, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h346, 12'h346, 12'h346, 12'h346, 12'h356, 12'h346, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h346, 12'h346, 12'h456, 12'h556, 12'h556, 12'h455, 12'h455, 12'h445, 12'h345, 12'h344, 12'h234, 12'h234, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h556, 12'h556, 12'h466, 12'h457, 12'h567, 12'h567, 12'h457, 12'h457, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h678, 12'h778, 12'h788, 12'h889, 12'h899, 12'h9aa, 12'haab, 12'hbbb, 12'hccc, 12'hcdd, 12'hddd, 
12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hbcd, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h99c, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'habc, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hbcd, 12'habc, 12'haab, 12'h9ab, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'h99b, 12'h99c, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'h9ab, 12'haab, 12'habc, 12'hbbc, 12'hbcc, 12'hccc, 12'hccc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hcdd, 12'hbbb, 12'h99a, 12'h89a, 12'h9ab, 12'h9ab, 12'h89a, 12'h78a, 12'h78a, 12'h78b, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h78c, 12'h78c, 12'h78c, 12'h78c, 12'h78c, 12'h78c, 12'h88d, 12'h88d, 12'h89d, 12'h99e, 12'h9ae, 
12'h9af, 12'habf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h9ae, 12'h8ae, 12'h8ae, 12'h8ae, 12'h7ae, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8bd, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'habd, 12'hbce, 12'hcdf, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heef, 12'hdef, 
12'hdde, 12'hcde, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h79b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hccc, 12'hbcc, 12'hbbb, 12'haaa, 12'h99a, 12'h899, 12'h888, 12'h778, 12'h677, 12'h567, 12'h566, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h345, 12'h345, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h245, 12'h345, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h346, 12'h346, 12'h345, 12'h345, 12'h345, 12'h345, 12'h245, 12'h245, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h566, 12'h556, 12'h456, 12'h455, 12'h445, 12'h345, 12'h345, 12'h334, 12'h234, 12'h234, 12'h334, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h457, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h678, 12'h778, 12'h788, 12'h889, 12'h999, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 
12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hbcd, 12'hbbd, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'haac, 12'habc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hdde, 12'hccd, 12'habc, 12'haab, 12'h9ab, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h9ab, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'haab, 12'habc, 12'hbbc, 12'hbcc, 12'hccd, 12'hccd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbc, 12'haab, 12'haab, 12'haab, 12'h9aa, 12'h89a, 12'h689, 12'h78a, 12'h79b, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h78b, 12'h68b, 12'h78c, 12'h78c, 12'h78c, 12'h78c, 12'h78c, 12'h89d, 12'h89d, 12'h89d, 12'h99d, 12'h9ae, 12'h9ae, 12'h9ae, 
12'habf, 12'habf, 12'h9bf, 12'h9ae, 12'h8ae, 12'h8ae, 12'h8ad, 12'h7ad, 12'h8ad, 12'h8ae, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h9be, 12'h9be, 12'h9bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'habd, 12'hbce, 12'hddf, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heef, 12'heef, 
12'hdef, 12'hdde, 12'hcde, 12'hcce, 12'hbcd, 12'hbbd, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h8ac, 12'h9ad, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hccc, 12'hbbc, 12'hbbb, 12'haaa, 12'h999, 12'h889, 12'h778, 12'h677, 12'h667, 12'h567, 12'h566, 12'h556, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h445, 12'h345, 12'h245, 12'h245, 12'h235, 12'h235, 12'h245, 12'h245, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h346, 12'h346, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h356, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h455, 12'h445, 12'h345, 12'h344, 12'h234, 12'h234, 12'h234, 12'h234, 12'h345, 12'h345, 12'h455, 12'h456, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h566, 12'h556, 12'h556, 12'h556, 12'h456, 12'h566, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h678, 12'h778, 12'h788, 12'h889, 12'h99a, 12'haaa, 12'habb, 12'hbcc, 12'hccc, 
12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hcde, 12'hccd, 12'hbcd, 12'habc, 12'haac, 12'h9ac, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'hccd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdee, 12'hccd, 12'habc, 12'haab, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h89b, 12'h99b, 12'h89b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 
12'h99c, 12'h9ac, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'haac, 12'habc, 12'hbcc, 12'hccd, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'habb, 12'h89a, 12'h78a, 12'h89b, 12'h89b, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79c, 12'h79b, 12'h79b, 12'h79b, 12'h78b, 12'h68b, 12'h68b, 12'h68b, 12'h68c, 12'h78c, 12'h78c, 12'h79c, 12'h89d, 12'h89d, 12'h99d, 12'h99d, 12'h9ae, 12'h9ae, 12'haae, 12'habe, 
12'haae, 12'h9ae, 12'h9ae, 12'h8ae, 12'h8ae, 12'h8ad, 12'h7ad, 12'h7ad, 12'h8ad, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8ae, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h89d, 12'h89d, 12'h8ad, 12'h9ad, 12'habd, 12'hbce, 12'hdef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 
12'hdef, 12'hdef, 12'hdde, 12'hcde, 12'hcce, 12'hbcd, 12'habd, 12'habc, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h8ab, 12'h8ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h89c, 12'h89c, 12'h8ac, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bd, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcdd, 12'hcde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbcc, 12'habb, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h677, 12'h567, 12'h566, 12'h456, 12'h456, 12'h556, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h445, 12'h345, 12'h345, 12'h245, 12'h245, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h346, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h346, 12'h446, 12'h456, 12'h356, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h455, 12'h445, 12'h345, 12'h234, 12'h234, 12'h234, 12'h234, 12'h345, 12'h445, 12'h456, 12'h556, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h567, 12'h567, 12'h677, 12'h778, 12'h788, 12'h889, 12'h99a, 12'haaa, 12'hbbb, 12'hccc, 
12'hccd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heee, 12'heee, 12'hdde, 12'hdde, 12'hcde, 12'hccd, 12'hbbd, 12'habc, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'habc, 12'hccd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hcdd, 12'hbbc, 12'habb, 12'haab, 12'h9ab, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h89b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 
12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h88a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'haac, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbc, 12'h99a, 12'h89a, 12'h89b, 12'h8ab, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79b, 12'h68b, 12'h68b, 12'h68b, 12'h67b, 12'h67b, 12'h68b, 12'h68b, 12'h78c, 12'h79c, 12'h89d, 12'h89d, 12'h89d, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ae, 12'h9ae, 12'h9ae, 12'h9ae, 
12'h9ae, 12'h9ae, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 12'h8ad, 12'h8ad, 12'h8be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h9be, 12'h8be, 12'h9be, 12'h8be, 12'h8ad, 12'h8ad, 12'h8ad, 12'h89d, 12'h89d, 12'h89c, 12'h89d, 12'h9ad, 12'habd, 12'hcde, 12'hdef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 
12'heef, 12'hdef, 12'hdef, 12'hdde, 12'hcde, 12'hccd, 12'hbcd, 12'hbcd, 12'habd, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ab, 12'h9ac, 12'h8ab, 12'h8ab, 12'h8ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h89c, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h89c, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bd, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hdee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'hddd, 12'hccd, 12'hbcc, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h667, 12'h667, 12'h566, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h455, 12'h555, 12'h556, 12'h556, 12'h455, 12'h445, 12'h445, 12'h334, 12'h234, 12'h234, 12'h334, 12'h345, 12'h455, 12'h456, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h567, 12'h667, 12'h678, 12'h788, 12'h889, 12'h99a, 12'haaa, 12'hbbb, 
12'hccc, 12'hcdd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'hdde, 12'hdde, 12'hcdd, 12'hccd, 12'hbcd, 12'hbbc, 12'hbbc, 12'hbcd, 12'hccd, 12'hdee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccc, 12'hbbc, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 
12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h78a, 12'h88a, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'haab, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hcdd, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'habb, 12'h99a, 12'h89b, 12'h8ab, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79b, 12'h79b, 12'h68b, 12'h68b, 12'h68b, 12'h68b, 12'h68b, 12'h79c, 12'h79c, 12'h89d, 12'h89d, 12'h89d, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ae, 12'h9ad, 
12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h7ad, 12'h7ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h8ad, 12'h79d, 12'h79d, 12'h79c, 12'h89c, 12'h9ad, 12'hbce, 12'hddf, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'heff, 12'heef, 12'hdef, 12'hdef, 12'hdde, 12'hcde, 12'hcce, 12'hbcd, 12'hbcd, 12'habd, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h89c, 12'h9ac, 12'h9ac, 12'h89c, 12'h9ac, 12'h99c, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hcdd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h889, 12'h788, 12'h677, 12'h667, 12'h667, 12'h566, 12'h566, 12'h566, 12'h556, 12'h456, 12'h456, 12'h456, 12'h556, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h456, 12'h455, 12'h455, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h555, 12'h556, 12'h556, 12'h556, 12'h556, 12'h455, 12'h445, 12'h345, 12'h234, 12'h234, 12'h334, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h567, 12'h667, 12'h678, 12'h789, 12'h889, 12'h99a, 12'haab, 
12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heef, 12'heff, 12'heff, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'hcdd, 12'hbbc, 12'habc, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'haac, 12'habc, 12'hbbc, 12'hbbc, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haab, 12'h9ab, 12'h9ab, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79c, 12'h79c, 12'h79b, 12'h79b, 12'h78c, 12'h79c, 12'h79c, 12'h79c, 12'h89d, 12'h89d, 12'h89d, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 
12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h7ad, 12'h79d, 12'h79c, 12'h79c, 12'h89d, 12'habd, 12'hcde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heff, 12'heef, 12'hdef, 12'hdee, 12'hdde, 12'hcde, 12'hccd, 12'hbcd, 12'hbcd, 12'habd, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h9ac, 12'h8ac, 12'h89c, 12'h8ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'habd, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'habb, 12'h9aa, 12'h899, 12'h888, 12'h788, 12'h778, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h566, 12'h556, 12'h556, 12'h456, 12'h455, 12'h445, 12'h345, 12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h345, 12'h345, 12'h445, 12'h445, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h555, 12'h555, 12'h556, 12'h556, 12'h566, 12'h566, 12'h556, 12'h556, 12'h455, 12'h345, 12'h345, 12'h334, 12'h234, 12'h234, 12'h345, 12'h345, 12'h345, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h677, 12'h778, 12'h789, 12'h899, 12'haaa, 
12'habb, 12'hbcc, 12'hccd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccd, 12'hbbc, 12'habb, 12'haab, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ac, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbcc, 12'habb, 12'haab, 12'h9bc, 12'h9bc, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89d, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 
12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h79d, 12'h79c, 12'h79c, 12'h79c, 12'h8ad, 12'hbce, 12'hdef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdef, 12'hdee, 12'hcde, 12'hcde, 12'hccd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89c, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habc, 12'habd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbce, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdee, 12'hdee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h899, 12'h888, 12'h788, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h677, 12'h667, 12'h666, 12'h566, 12'h556, 12'h555, 12'h445, 12'h445, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h455, 12'h445, 12'h345, 12'h455, 12'h455, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h566, 12'h566, 12'h666, 12'h566, 12'h566, 12'h556, 12'h455, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h567, 12'h667, 12'h678, 12'h788, 12'h889, 12'h99a, 
12'haab, 12'hbbb, 12'hccc, 12'hcdd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccd, 12'hbbc, 12'habb, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89a, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ac, 12'haac, 12'habc, 12'hbbd, 12'hccd, 12'hccd, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hccc, 12'hbbc, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h89c, 
12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h7ad, 12'h8ad, 12'h79d, 12'h79c, 12'h79c, 12'h89c, 12'habd, 12'hcde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdef, 12'hdee, 12'hdde, 12'hcde, 12'hcce, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'habd, 12'habd, 12'h9bc, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'habc, 12'habd, 12'hacd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdee, 12'hdee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h777, 12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h566, 12'h566, 12'h566, 12'h556, 12'h566, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h555, 12'h555, 12'h555, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 
12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h456, 12'h455, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h555, 12'h555, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h456, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h567, 12'h567, 12'h668, 12'h778, 12'h789, 12'h899, 
12'h9aa, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'hccc, 12'hbbc, 12'haab, 12'h9ab, 12'h99b, 12'h99b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h99b, 12'h99b, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'haac, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hcde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbcc, 12'habc, 12'habc, 12'h9bc, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 
12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h8ad, 12'h8ad, 12'h8ae, 12'h8be, 12'h8be, 12'h8be, 12'h8bf, 12'h8bf, 12'h8be, 12'h8bf, 12'h8bf, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h7ad, 12'h7ad, 12'h79d, 12'h79c, 12'h79c, 12'h9ad, 12'hbce, 12'hdef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hcde, 12'hccd, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'habd, 12'habd, 12'habd, 12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'habc, 12'habd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h666, 12'h556, 12'h445, 12'h455, 12'h445, 12'h444, 12'h444, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h555, 12'h555, 12'h556, 12'h566, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h677, 12'h677, 12'h677, 12'h777, 12'h777, 12'h778, 12'h778, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 
12'h566, 12'h566, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h455, 12'h455, 12'h555, 12'h555, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h455, 12'h455, 12'h445, 12'h345, 12'h445, 12'h455, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h557, 12'h567, 12'h667, 12'h678, 12'h778, 12'h889, 
12'h99a, 12'haaa, 12'hbbb, 12'hccc, 12'hccd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'habc, 12'haab, 12'h9ab, 12'h99b, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'haac, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbbc, 12'habc, 12'h9bc, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 
12'h89c, 12'h89c, 12'h79c, 12'h89d, 12'h8ad, 12'h8ae, 12'h9be, 12'h9bf, 12'h9bf, 12'h9bf, 12'h8bf, 12'h8bf, 12'h8cf, 12'h8bf, 12'h8bf, 12'h8bf, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h7ad, 12'h79d, 12'h79c, 12'h79c, 12'h89c, 12'haad, 12'hcde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hcde, 12'hcde, 12'hbcd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habc, 12'habc, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdee, 12'hdee, 12'heee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'h566, 12'h455, 12'h344, 12'h233, 12'h233, 12'h223, 12'h223, 12'h223, 12'h223, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h333, 12'h334, 12'h344, 12'h344, 12'h445, 12'h455, 12'h555, 12'h555, 12'h556, 12'h566, 12'h566, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h677, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h677, 
12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h456, 12'h455, 12'h455, 12'h455, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h555, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h456, 12'h445, 12'h445, 12'h345, 12'h344, 12'h345, 12'h455, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h557, 12'h567, 12'h667, 12'h678, 12'h789, 
12'h889, 12'h99a, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbbc, 12'haab, 12'haab, 12'h99b, 12'h99a, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'haac, 12'haac, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccd, 12'hbbc, 12'habc, 12'h9bc, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 12'h89c, 12'h89c, 12'h89c, 12'h89c, 12'h79c, 12'h79c, 12'h79c, 
12'h89c, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ae, 12'h9be, 12'h9bf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9bf, 12'h8bf, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h7ad, 12'h79d, 12'h79c, 12'h79c, 12'h9ad, 12'hbce, 12'hdef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hcde, 12'hcde, 12'hccd, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'habc, 12'habc, 12'hbbd, 12'hbcd, 12'hccd, 12'hccd, 12'hcde, 12'hcde, 12'hdde, 12'hdee, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h666, 12'h445, 12'h334, 12'h233, 12'h223, 12'h122, 12'h112, 12'h122, 12'h112, 12'h122, 12'h122, 12'h122, 12'h123, 12'h223, 12'h223, 12'h233, 12'h233, 12'h233, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h344, 12'h344, 12'h334, 12'h334, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h444, 12'h344, 12'h344, 12'h334, 12'h344, 12'h444, 12'h444, 12'h455, 12'h555, 12'h555, 12'h556, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h778, 
12'h778, 12'h778, 12'h778, 12'h778, 12'h788, 12'h788, 12'h778, 12'h778, 12'h677, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h455, 12'h455, 12'h455, 12'h555, 12'h555, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h456, 12'h455, 12'h445, 12'h345, 12'h345, 12'h455, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h567, 12'h567, 12'h668, 12'h778, 
12'h889, 12'h99a, 12'haaa, 12'hbbb, 12'hbcc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'haab, 12'h9ab, 12'h99a, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'habc, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hccd, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'hbcc, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h89c, 12'h79c, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 
12'h8ad, 12'h8ad, 12'h8ad, 12'h9ae, 12'h9be, 12'h9be, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ad, 12'h8ad, 12'h79d, 12'h79c, 12'h89c, 12'habd, 12'hdde, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdef, 12'hdee, 12'hdde, 12'hcde, 12'hcde, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h9ab, 12'haac, 12'habc, 12'habc, 12'hbbd, 12'hbcd, 12'hccd, 12'hcdd, 12'hcde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h777, 12'h666, 12'h555, 12'h444, 12'h333, 12'h222, 12'h122, 12'h112, 12'h112, 12'h112, 12'h112, 12'h111, 12'h111, 12'h112, 12'h112, 12'h122, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h122, 12'h112, 12'h011, 12'h011, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h122, 12'h222, 12'h222, 12'h222, 12'h223, 12'h333, 12'h333, 12'h444, 12'h444, 12'h444, 12'h555, 12'h555, 12'h555, 12'h555, 12'h556, 12'h566, 12'h666, 12'h666, 12'h566, 12'h666, 12'h566, 12'h666, 12'h666, 12'h667, 12'h667, 12'h667, 12'h667, 
12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h667, 12'h666, 12'h566, 12'h566, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h557, 12'h557, 12'h567, 12'h678, 
12'h778, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'hbbb, 12'haab, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h89b, 12'h99b, 
12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'haac, 12'habc, 12'habc, 12'hbbc, 12'hbbd, 12'hbcd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'hbbc, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 
12'h8ad, 12'h8ad, 12'h8ad, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9bf, 12'h9bf, 12'h9bf, 12'h8bf, 12'h8be, 12'h8be, 12'h8be, 12'h8ae, 12'h8ad, 12'h8ad, 12'h89c, 12'h89c, 12'haad, 12'hcce, 12'hdef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'hdef, 12'hdee, 12'hdde, 12'hcde, 12'hccd, 12'hbcd, 12'hbcd, 12'habc, 12'habc, 12'habc, 12'habc, 12'haac, 12'h9ab, 12'h9ab, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbcd, 12'hbcd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h555, 12'h444, 12'h333, 12'h222, 12'h222, 12'h122, 12'h111, 12'h112, 12'h112, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h112, 12'h122, 12'h122, 12'h122, 12'h121, 12'h121, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h001, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 
12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h555, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h666, 12'h666, 12'h667, 12'h667, 12'h677, 12'h777, 12'h777, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h788, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h788, 12'h788, 12'h778, 12'h778, 12'h777, 12'h677, 12'h667, 12'h667, 12'h566, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h556, 12'h556, 12'h566, 12'h566, 12'h567, 12'h567, 12'h567, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h566, 12'h566, 12'h466, 12'h467, 12'h467, 12'h467, 12'h467, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h567, 12'h667, 
12'h678, 12'h788, 12'h899, 12'h9aa, 12'habb, 12'hbcc, 12'hcdd, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hddd, 12'hbbb, 12'h9aa, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ab, 
12'h9ab, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'habc, 12'hbbc, 12'hbbd, 12'hbcd, 12'hccd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hcdd, 12'hbcd, 12'habc, 12'habc, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h8ad, 
12'h8ad, 12'h8ad, 12'h8ad, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9ce, 12'h9ce, 12'h9cf, 12'h9cf, 12'h9cf, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h9ad, 12'hbce, 12'hdee, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hcde, 12'hcde, 12'hcde, 12'hbcd, 12'hbbd, 12'habc, 12'habc, 12'haac, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'haac, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hbcd, 12'hccd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccb, 12'haaa, 12'h999, 12'h777, 12'h666, 12'h555, 12'h444, 12'h333, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h101, 12'h101, 12'h000, 12'h000, 12'h001, 12'h001, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h222, 12'h333, 12'h333, 12'h333, 12'h333, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h001, 12'h002, 12'h002, 12'h002, 12'h002, 12'h002, 12'h012, 12'h012, 12'h012, 
12'h022, 12'h023, 12'h023, 12'h123, 12'h123, 12'h123, 12'h223, 12'h334, 12'h445, 12'h445, 12'h445, 12'h445, 12'h455, 12'h455, 12'h555, 12'h556, 12'h556, 12'h566, 12'h666, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h677, 12'h677, 12'h677, 12'h667, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h667, 12'h667, 12'h667, 12'h677, 12'h677, 12'h678, 12'h678, 12'h678, 12'h678, 12'h678, 12'h677, 12'h677, 12'h677, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h457, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h557, 12'h567, 
12'h667, 12'h678, 12'h889, 12'h99a, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdde, 12'hbbc, 12'h9aa, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ab, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 
12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbd, 12'hbcd, 12'hccd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hdde, 12'hccd, 12'hbcd, 12'habc, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8bd, 12'h9bd, 12'h9ad, 12'h9ad, 
12'h8ad, 12'h8ad, 12'h8bd, 12'h8be, 12'h9be, 12'h9be, 12'h8be, 12'h9ce, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8be, 12'h8bd, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'hbcd, 12'hdde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'hdee, 12'hdee, 12'hdde, 12'hcde, 12'hcdd, 12'hbcd, 12'hbcd, 12'habc, 12'habc, 12'haab, 12'haab, 12'haab, 12'habb, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbcc, 12'hbcd, 12'hccd, 12'hcdd, 12'hddd, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'h555, 12'h444, 12'h333, 12'h232, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h023, 12'h123, 
12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h233, 12'h234, 12'h234, 12'h234, 12'h234, 12'h233, 12'h333, 12'h334, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h344, 12'h444, 12'h444, 12'h444, 12'h444, 12'h344, 12'h344, 12'h345, 12'h445, 12'h455, 12'h455, 12'h556, 12'h556, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h667, 12'h667, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h778, 12'h778, 12'h778, 12'h788, 12'h788, 12'h788, 12'h788, 12'h788, 12'h778, 12'h778, 12'h778, 12'h678, 12'h677, 12'h677, 12'h677, 12'h677, 12'h677, 12'h667, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h557, 12'h557, 12'h457, 12'h557, 12'h557, 12'h567, 
12'h667, 12'h677, 12'h788, 12'h899, 12'h9aa, 12'hbbb, 12'hccc, 12'hcdd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccd, 12'haab, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89b, 12'h89b, 12'h89a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'haac, 12'habc, 12'habc, 12'habc, 12'hbbc, 
12'hbbc, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdde, 12'hccd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h9bd, 12'h9bd, 12'h8ad, 
12'h8ad, 12'h8ad, 12'h8bd, 12'h8be, 12'h9be, 12'h9be, 12'h8be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h9be, 12'h8be, 12'h8be, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'hbcd, 12'hdde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hcde, 12'hcdd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hbcc, 12'hccd, 12'hccd, 12'hcdd, 12'hddd, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h666, 12'h554, 12'h343, 12'h333, 12'h222, 12'h221, 12'h121, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h211, 12'h211, 12'h221, 12'h222, 12'h211, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h023, 12'h123, 12'h123, 12'h123, 
12'h123, 12'h012, 12'h112, 12'h112, 12'h112, 12'h012, 12'h012, 12'h022, 12'h123, 12'h123, 12'h112, 12'h112, 12'h112, 12'h112, 12'h112, 12'h112, 12'h122, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h122, 12'h112, 12'h012, 12'h012, 12'h012, 12'h122, 12'h123, 12'h123, 12'h233, 12'h334, 12'h344, 12'h444, 12'h445, 12'h445, 12'h455, 12'h455, 12'h455, 12'h456, 12'h556, 12'h566, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h667, 12'h677, 12'h778, 12'h778, 
12'h778, 12'h778, 12'h888, 12'h999, 12'haaa, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'hdee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hccc, 12'haab, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ac, 12'haab, 12'haac, 12'haac, 12'haac, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 
12'hccd, 12'hcdd, 12'hcdd, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hcde, 12'hccd, 12'hbcd, 12'habd, 12'habd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 
12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9be, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9ad, 12'habd, 12'hbcd, 12'hdde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heff, 12'heef, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hcdd, 12'hcdd, 12'hccd, 12'hccd, 12'hccd, 12'hcdd, 12'hcdd, 12'hddd, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h888, 12'h777, 12'h555, 12'h444, 12'h233, 12'h222, 12'h222, 12'h222, 12'h122, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h221, 12'h221, 12'h221, 12'h211, 12'h211, 12'h211, 12'h211, 12'h211, 12'h221, 12'h221, 12'h221, 12'h221, 12'h221, 12'h221, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h222, 12'h222, 12'h223, 
12'h223, 12'h212, 12'h212, 12'h212, 12'h112, 12'h112, 12'h112, 12'h112, 12'h222, 12'h212, 12'h212, 12'h111, 12'h102, 12'h102, 12'h112, 12'h222, 12'h222, 12'h222, 12'h112, 12'h112, 12'h111, 12'h101, 12'h111, 12'h112, 12'h222, 12'h222, 12'h122, 12'h121, 12'h122, 12'h122, 12'h122, 12'h122, 12'h222, 12'h223, 12'h233, 12'h233, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h445, 12'h344, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h335, 12'h335, 12'h334, 12'h335, 12'h345, 12'h445, 12'h445, 12'h445, 12'h555, 12'h555, 12'h556, 12'h656, 12'h666, 12'h666, 12'h666, 12'h667, 12'h667, 12'h767, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h878, 12'h888, 
12'h888, 12'h888, 12'h888, 12'h999, 12'h99a, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hddd, 12'hbbc, 12'h99a, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'habb, 12'habc, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcdd, 12'hddd, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdde, 12'hcde, 12'hcce, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ad, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 
12'h8ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h8bd, 12'h8bd, 12'h8bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'hcde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h777, 12'h666, 12'h455, 12'h334, 12'h233, 12'h223, 12'h112, 12'h112, 12'h112, 12'h222, 12'h222, 12'h222, 12'h122, 12'h111, 12'h111, 12'h111, 12'h111, 12'h112, 12'h111, 12'h111, 12'h111, 12'h111, 12'h011, 12'h011, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h211, 12'h221, 12'h221, 12'h222, 12'h222, 12'h221, 12'h221, 12'h221, 12'h221, 12'h221, 12'h211, 12'h211, 12'h211, 12'h211, 12'h321, 12'h321, 12'h321, 12'h320, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h322, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h312, 12'h312, 12'h312, 12'h322, 12'h323, 
12'h323, 12'h323, 12'h322, 12'h212, 12'h212, 12'h211, 12'h211, 12'h212, 12'h322, 12'h222, 12'h212, 12'h211, 12'h212, 12'h212, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h212, 12'h212, 12'h211, 12'h212, 12'h222, 12'h333, 12'h333, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h122, 12'h222, 12'h222, 12'h222, 12'h222, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h113, 12'h113, 12'h113, 12'h223, 12'h223, 12'h223, 12'h224, 12'h224, 12'h224, 12'h113, 12'h113, 12'h224, 12'h224, 12'h334, 12'h335, 12'h444, 12'h444, 12'h445, 12'h545, 12'h555, 12'h555, 12'h556, 12'h656, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h667, 12'h767, 12'h777, 
12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'hdde, 12'hcdd, 12'habb, 12'habb, 12'habb, 12'haab, 12'habb, 12'habb, 12'habc, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcdd, 12'hcdd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hdde, 12'hcde, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'h9bd, 12'h9ac, 12'h9ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 
12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ad, 12'h8ad, 12'h9ad, 12'h9ad, 12'h9bd, 12'h9ad, 12'h9ad, 12'h9ad, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'hcde, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heff, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h667, 12'h556, 12'h445, 12'h334, 12'h223, 12'h113, 12'h002, 12'h002, 12'h012, 12'h122, 12'h222, 12'h222, 12'h122, 12'h111, 12'h011, 12'h111, 12'h111, 12'h112, 12'h122, 12'h122, 12'h112, 12'h112, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h211, 12'h221, 12'h222, 12'h222, 12'h222, 12'h222, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h321, 12'h322, 12'h323, 12'h323, 12'h312, 12'h312, 12'h312, 12'h212, 12'h312, 12'h312, 12'h312, 12'h323, 
12'h323, 12'h323, 12'h322, 12'h322, 12'h222, 12'h222, 12'h222, 12'h212, 12'h222, 12'h222, 12'h212, 12'h211, 12'h212, 12'h212, 12'h222, 12'h322, 12'h323, 12'h323, 12'h333, 12'h323, 12'h323, 12'h333, 12'h333, 12'h333, 12'h444, 12'h434, 12'h333, 12'h232, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h233, 12'h233, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h233, 12'h223, 12'h223, 12'h223, 12'h113, 12'h002, 12'h002, 12'h002, 12'h112, 12'h223, 12'h223, 12'h224, 12'h224, 12'h224, 12'h223, 12'h113, 12'h113, 12'h103, 12'h113, 12'h214, 12'h223, 12'h223, 12'h322, 12'h323, 12'h333, 12'h333, 12'h333, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h444, 12'h444, 12'h444, 12'h444, 
12'h444, 12'h545, 12'h555, 12'h666, 12'h666, 12'h878, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'heee, 12'hdde, 12'hccc, 12'hbcc, 12'hbcc, 12'hbbc, 12'hbcc, 12'hbcc, 12'hbcc, 12'hbcc, 12'hbcc, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcdd, 12'hcdd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 
12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hdde, 12'hcce, 12'hbcd, 12'habd, 12'habd, 12'h9ad, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ad, 12'h8ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ad, 
12'h9ad, 12'h9ad, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9bd, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'hcde, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccd, 12'hbbb, 12'haaa, 12'h999, 12'h778, 12'h666, 12'h556, 12'h445, 12'h334, 12'h223, 12'h112, 12'h002, 12'h002, 12'h002, 12'h112, 12'h112, 12'h112, 12'h111, 12'h011, 12'h011, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h112, 12'h212, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h321, 12'h321, 12'h321, 12'h322, 12'h322, 12'h332, 12'h332, 12'h332, 12'h332, 12'h322, 12'h312, 12'h212, 12'h202, 12'h212, 12'h212, 12'h202, 12'h212, 12'h212, 12'h312, 12'h323, 
12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h322, 12'h222, 12'h222, 12'h222, 12'h212, 12'h222, 12'h222, 12'h322, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h434, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h333, 12'h232, 12'h232, 12'h222, 12'h222, 12'h222, 12'h233, 12'h233, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h223, 12'h223, 12'h112, 12'h002, 12'h002, 12'h113, 12'h113, 12'h223, 12'h334, 12'h334, 12'h334, 12'h334, 12'h224, 12'h223, 12'h213, 12'h113, 12'h113, 12'h213, 12'h213, 12'h112, 12'h211, 12'h212, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h212, 12'h211, 12'h211, 12'h211, 12'h211, 12'h222, 12'h222, 12'h222, 12'h322, 
12'h222, 12'h322, 12'h333, 12'h444, 12'h555, 12'h666, 12'h777, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heee, 12'hddd, 12'hcdd, 12'hcdd, 12'hcdd, 12'hcdd, 12'hcdd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'heff, 
12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdde, 12'hcde, 12'hbcd, 12'habd, 12'habd, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h8ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 
12'h9ad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'habd, 12'hbcd, 12'hcde, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h556, 12'h555, 12'h445, 12'h334, 12'h223, 12'h012, 12'h002, 12'h002, 12'h012, 12'h002, 12'h001, 12'h011, 12'h012, 12'h012, 12'h011, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h332, 12'h332, 12'h322, 12'h322, 12'h322, 12'h212, 12'h202, 12'h202, 12'h202, 12'h202, 12'h202, 12'h212, 12'h212, 12'h212, 12'h212, 
12'h212, 12'h212, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h232, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h233, 12'h223, 12'h223, 12'h223, 12'h222, 12'h222, 12'h222, 12'h222, 12'h223, 12'h223, 12'h223, 12'h112, 12'h213, 12'h113, 12'h223, 12'h223, 12'h223, 12'h323, 12'h323, 12'h223, 12'h213, 12'h213, 12'h213, 12'h213, 12'h223, 12'h223, 12'h223, 12'h222, 12'h222, 12'h332, 12'h332, 12'h333, 12'h332, 12'h332, 12'h322, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h322, 12'h333, 12'h333, 
12'h222, 12'h222, 12'h333, 12'h444, 12'h544, 12'h555, 12'h777, 12'h888, 12'h999, 12'haaa, 12'hccc, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hcde, 12'hbcd, 12'habd, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ad, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 
12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bd, 12'habd, 12'hbbd, 12'hbcd, 12'hcde, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'haab, 12'h999, 12'h888, 12'h667, 12'h555, 12'h445, 12'h334, 12'h223, 12'h123, 12'h002, 12'h112, 12'h123, 12'h123, 12'h112, 12'h002, 12'h112, 12'h122, 12'h122, 12'h112, 12'h122, 12'h122, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h322, 12'h212, 12'h212, 12'h212, 12'h212, 12'h202, 12'h212, 12'h212, 12'h212, 12'h202, 12'h211, 
12'h211, 12'h211, 12'h211, 12'h211, 12'h212, 12'h212, 12'h212, 12'h222, 12'h222, 12'h323, 12'h323, 12'h323, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h122, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h111, 12'h111, 12'h112, 12'h122, 12'h222, 12'h212, 12'h212, 12'h112, 12'h111, 12'h111, 12'h111, 12'h112, 12'h223, 12'h323, 12'h223, 12'h223, 12'h222, 12'h222, 12'h222, 12'h223, 12'h223, 12'h223, 12'h223, 12'h213, 12'h213, 12'h223, 12'h223, 12'h223, 12'h323, 12'h333, 12'h333, 12'h332, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h332, 12'h232, 12'h222, 12'h222, 12'h222, 12'h232, 12'h332, 12'h333, 12'h333, 12'h333, 
12'h222, 12'h221, 12'h222, 12'h333, 12'h444, 12'h555, 12'h666, 12'h787, 12'h898, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hcde, 12'hbcd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h8ac, 12'h9ac, 
12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'hbbd, 12'hbcd, 12'hcde, 12'hdee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hbbb, 12'haaa, 12'h999, 12'h777, 12'h666, 12'h455, 12'h334, 12'h224, 12'h113, 12'h113, 12'h002, 12'h223, 12'h233, 12'h334, 12'h223, 12'h122, 12'h223, 12'h333, 12'h233, 12'h123, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h022, 12'h122, 12'h112, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h222, 12'h222, 12'h112, 12'h112, 12'h112, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h322, 12'h322, 12'h322, 12'h322, 12'h222, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h102, 12'h102, 12'h101, 
12'h101, 12'h101, 12'h101, 12'h111, 12'h111, 12'h111, 12'h112, 12'h222, 12'h222, 12'h223, 12'h223, 12'h223, 12'h222, 12'h222, 12'h222, 12'h122, 12'h112, 12'h112, 12'h122, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h122, 12'h122, 12'h222, 12'h232, 12'h222, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h122, 12'h222, 12'h122, 12'h112, 12'h112, 12'h112, 12'h111, 12'h111, 12'h112, 12'h222, 12'h323, 12'h333, 12'h333, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h323, 12'h323, 12'h333, 12'h334, 12'h334, 12'h333, 12'h232, 12'h332, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h222, 12'h232, 12'h232, 12'h232, 12'h232, 12'h332, 12'h333, 12'h333, 12'h333, 
12'h232, 12'h232, 12'h232, 12'h333, 12'h444, 12'h454, 12'h665, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hccc, 12'hddc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hcde, 12'hbcd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h9ac, 12'h9ac, 
12'h9bc, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbcd, 12'hcde, 12'hdee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h556, 12'h445, 12'h334, 12'h223, 12'h223, 12'h223, 12'h223, 12'h334, 12'h445, 12'h555, 12'h445, 12'h445, 12'h445, 12'h556, 12'h455, 12'h445, 12'h344, 12'h334, 12'h233, 12'h223, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h122, 12'h112, 12'h112, 12'h112, 12'h112, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h212, 12'h213, 12'h213, 12'h223, 12'h213, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h212, 12'h112, 12'h112, 12'h112, 
12'h101, 12'h101, 12'h101, 12'h101, 12'h112, 12'h112, 12'h112, 12'h112, 12'h112, 12'h112, 12'h122, 12'h223, 12'h122, 12'h222, 12'h222, 12'h122, 12'h122, 12'h122, 12'h223, 12'h233, 12'h333, 12'h333, 12'h333, 12'h333, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h223, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h333, 12'h333, 12'h334, 12'h333, 12'h232, 12'h232, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h232, 12'h232, 12'h232, 12'h232, 12'h332, 12'h332, 12'h333, 12'h333, 
12'h332, 12'h232, 12'h232, 12'h333, 12'h443, 12'h454, 12'h565, 12'h676, 12'h887, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'hdee, 12'hdde, 12'hccd, 12'hbbd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 12'h9bc, 
12'habc, 12'habc, 12'habc, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hccd, 12'hdde, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h888, 12'h667, 12'h455, 12'h344, 12'h334, 12'h234, 12'h334, 12'h334, 12'h334, 12'h455, 12'h667, 12'h677, 12'h667, 12'h667, 12'h677, 12'h778, 12'h677, 12'h666, 12'h555, 12'h445, 12'h344, 12'h234, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h123, 12'h123, 12'h123, 12'h123, 12'h223, 12'h223, 12'h123, 12'h123, 12'h223, 12'h123, 12'h223, 12'h223, 12'h123, 12'h113, 12'h113, 12'h213, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h213, 12'h213, 12'h213, 12'h213, 12'h213, 12'h213, 12'h213, 12'h213, 12'h213, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h113, 12'h112, 12'h112, 
12'h112, 12'h112, 12'h112, 12'h112, 12'h012, 12'h112, 12'h112, 12'h112, 12'h012, 12'h012, 12'h122, 12'h123, 12'h123, 12'h223, 12'h122, 12'h022, 12'h122, 12'h122, 12'h223, 12'h233, 12'h333, 12'h333, 12'h333, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h223, 12'h222, 12'h222, 12'h222, 12'h223, 12'h233, 12'h333, 12'h333, 12'h333, 12'h333, 12'h223, 12'h223, 12'h222, 12'h223, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h232, 12'h232, 12'h222, 12'h221, 12'h221, 12'h221, 12'h221, 12'h221, 12'h221, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h332, 
12'h232, 12'h232, 12'h232, 12'h332, 12'h343, 12'h444, 12'h555, 12'h666, 12'h777, 12'h888, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heef, 12'heef, 12'hdde, 12'hcde, 12'hbcd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'habd, 12'habd, 12'habc, 12'habd, 12'habd, 
12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hcde, 12'hdde, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h888, 12'h666, 12'h445, 12'h344, 12'h334, 12'h334, 12'h334, 12'h345, 12'h445, 12'h556, 12'h777, 12'h888, 12'h788, 12'h788, 12'h888, 12'h889, 12'h888, 12'h777, 12'h566, 12'h455, 12'h445, 12'h334, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h234, 12'h234, 12'h234, 12'h234, 12'h334, 12'h334, 12'h234, 12'h223, 12'h223, 12'h223, 12'h224, 12'h334, 12'h334, 12'h334, 12'h234, 12'h224, 12'h224, 12'h224, 12'h224, 12'h214, 12'h214, 12'h224, 12'h224, 12'h224, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h123, 12'h123, 12'h123, 
12'h113, 12'h113, 12'h113, 12'h113, 12'h123, 12'h123, 12'h123, 12'h123, 12'h012, 12'h012, 12'h123, 12'h123, 12'h223, 12'h223, 12'h122, 12'h022, 12'h122, 12'h122, 12'h122, 12'h123, 12'h233, 12'h233, 12'h233, 12'h223, 12'h122, 12'h122, 12'h122, 12'h112, 12'h122, 12'h123, 12'h123, 12'h223, 12'h223, 12'h223, 12'h223, 12'h122, 12'h122, 12'h122, 12'h122, 12'h223, 12'h233, 12'h334, 12'h334, 12'h334, 12'h223, 12'h112, 12'h112, 12'h112, 12'h212, 12'h212, 12'h222, 12'h322, 12'h323, 12'h323, 12'h323, 12'h322, 12'h322, 12'h222, 12'h212, 12'h212, 12'h212, 12'h222, 12'h222, 12'h232, 12'h232, 12'h232, 12'h232, 12'h231, 12'h231, 12'h231, 12'h231, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 
12'h232, 12'h231, 12'h232, 12'h232, 12'h232, 12'h343, 12'h454, 12'h555, 12'h676, 12'h888, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'hdee, 12'hdde, 12'hcde, 12'hcde, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 
12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h999, 12'h777, 12'h556, 12'h444, 12'h344, 12'h334, 12'h334, 12'h345, 12'h445, 12'h455, 12'h667, 12'h788, 12'h899, 12'h899, 12'h899, 12'h99a, 12'h99a, 12'h899, 12'h788, 12'h667, 12'h556, 12'h445, 12'h345, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h345, 12'h335, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h334, 12'h234, 12'h224, 12'h224, 12'h224, 12'h224, 12'h224, 12'h224, 12'h224, 12'h124, 12'h123, 12'h123, 12'h124, 12'h224, 12'h223, 12'h224, 12'h224, 12'h224, 12'h224, 
12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h123, 12'h223, 12'h123, 12'h123, 12'h123, 12'h123, 12'h223, 12'h233, 12'h233, 12'h123, 12'h123, 12'h022, 12'h112, 12'h012, 12'h012, 12'h022, 12'h022, 12'h022, 12'h022, 12'h122, 12'h112, 12'h012, 12'h112, 12'h012, 12'h013, 12'h023, 12'h123, 12'h123, 12'h123, 12'h123, 12'h022, 12'h012, 12'h012, 12'h122, 12'h123, 12'h223, 12'h233, 12'h333, 12'h333, 12'h223, 12'h112, 12'h112, 12'h112, 12'h212, 12'h222, 12'h222, 12'h222, 12'h223, 12'h223, 12'h223, 12'h222, 12'h222, 12'h222, 12'h222, 12'h212, 12'h212, 12'h222, 12'h222, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 
12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h343, 12'h444, 12'h555, 12'h666, 12'h777, 12'h898, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddc, 12'hbbb, 12'haa9, 12'h888, 12'h667, 12'h455, 12'h344, 12'h334, 12'h334, 12'h334, 12'h345, 12'h455, 12'h556, 12'h667, 12'h788, 12'h999, 12'h99a, 12'h9aa, 12'h9aa, 12'h9aa, 12'h999, 12'h788, 12'h667, 12'h556, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h335, 12'h335, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h335, 12'h335, 12'h335, 12'h235, 12'h235, 12'h235, 12'h235, 12'h335, 12'h235, 12'h234, 12'h224, 12'h224, 12'h234, 12'h234, 12'h224, 12'h234, 12'h234, 12'h234, 12'h234, 
12'h224, 12'h224, 12'h224, 12'h124, 12'h124, 12'h123, 12'h123, 12'h123, 12'h223, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h123, 12'h123, 12'h023, 12'h012, 12'h012, 12'h013, 12'h023, 12'h023, 12'h123, 12'h234, 12'h234, 12'h234, 12'h124, 12'h124, 12'h023, 12'h023, 12'h023, 12'h023, 12'h123, 12'h123, 12'h013, 12'h012, 12'h112, 12'h112, 12'h112, 12'h113, 12'h223, 12'h223, 12'h223, 12'h233, 12'h233, 12'h234, 12'h334, 12'h233, 12'h323, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h323, 12'h323, 12'h333, 12'h323, 12'h323, 12'h323, 12'h232, 12'h232, 12'h232, 12'h232, 12'h232, 12'h132, 12'h232, 12'h232, 12'h232, 12'h232, 12'h233, 12'h333, 12'h333, 12'h333, 12'h233, 12'h232, 12'h232, 12'h232, 
12'h232, 12'h232, 12'h232, 12'h233, 12'h333, 12'h343, 12'h444, 12'h455, 12'h566, 12'h777, 12'h888, 12'h999, 12'haba, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hccc, 12'hbaa, 12'h999, 12'h777, 12'h666, 12'h445, 12'h334, 12'h334, 12'h234, 12'h234, 12'h345, 12'h445, 12'h456, 12'h667, 12'h778, 12'h889, 12'h99a, 12'h9aa, 12'haaa, 12'h9aa, 12'h899, 12'h788, 12'h667, 12'h556, 12'h445, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h335, 12'h335, 12'h335, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h446, 12'h446, 12'h446, 12'h446, 12'h345, 12'h345, 12'h445, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h346, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h235, 12'h235, 12'h235, 12'h335, 12'h335, 12'h235, 
12'h235, 12'h235, 12'h234, 12'h124, 12'h124, 12'h114, 12'h114, 12'h124, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h234, 12'h134, 12'h124, 12'h023, 12'h013, 12'h113, 12'h013, 12'h123, 12'h124, 12'h234, 12'h345, 12'h345, 12'h235, 12'h234, 12'h134, 12'h134, 12'h134, 12'h134, 12'h124, 12'h123, 12'h123, 12'h113, 12'h113, 12'h113, 12'h113, 12'h113, 12'h113, 12'h113, 12'h113, 12'h223, 12'h334, 12'h334, 12'h344, 12'h344, 12'h334, 12'h334, 12'h233, 12'h223, 12'h123, 12'h113, 12'h223, 12'h223, 12'h323, 12'h333, 12'h334, 12'h334, 12'h334, 12'h333, 12'h233, 12'h132, 12'h132, 12'h232, 12'h232, 12'h132, 12'h232, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h232, 12'h232, 12'h232, 
12'h232, 12'h232, 12'h232, 12'h233, 12'h233, 12'h333, 12'h344, 12'h454, 12'h555, 12'h666, 12'h788, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hedd, 12'hddc, 12'hcbb, 12'haaa, 12'h888, 12'h777, 12'h556, 12'h445, 12'h334, 12'h234, 12'h224, 12'h234, 12'h345, 12'h445, 12'h456, 12'h567, 12'h778, 12'h889, 12'h99a, 12'h9aa, 12'haab, 12'h9aa, 12'h899, 12'h778, 12'h567, 12'h456, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h335, 12'h335, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h446, 12'h456, 12'h456, 12'h456, 12'h446, 12'h346, 12'h346, 12'h446, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h446, 12'h446, 12'h346, 12'h446, 12'h446, 12'h346, 12'h346, 12'h346, 12'h446, 12'h446, 12'h446, 
12'h346, 12'h346, 12'h345, 12'h335, 12'h235, 12'h225, 12'h224, 12'h235, 12'h335, 12'h345, 12'h335, 12'h235, 12'h235, 12'h335, 12'h235, 12'h245, 12'h335, 12'h235, 12'h235, 12'h335, 12'h335, 12'h445, 12'h456, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h467, 12'h456, 12'h456, 12'h456, 12'h346, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h335, 12'h234, 12'h234, 12'h334, 12'h335, 12'h335, 12'h345, 12'h334, 12'h234, 12'h123, 12'h013, 12'h013, 12'h002, 12'h002, 12'h113, 12'h113, 12'h223, 12'h223, 12'h223, 12'h223, 12'h223, 12'h122, 12'h132, 12'h122, 12'h122, 12'h122, 12'h132, 12'h132, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h132, 12'h122, 12'h122, 12'h122, 
12'h122, 12'h122, 12'h122, 12'h123, 12'h122, 12'h233, 12'h343, 12'h344, 12'h455, 12'h566, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h777, 12'h666, 12'h555, 12'h444, 12'h344, 12'h334, 12'h234, 12'h334, 12'h445, 12'h556, 12'h556, 12'h667, 12'h778, 12'h789, 12'h99a, 12'haab, 12'haab, 12'h9aa, 12'h89a, 12'h778, 12'h567, 12'h456, 12'h446, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h335, 12'h335, 12'h235, 12'h335, 12'h335, 12'h345, 12'h345, 12'h346, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h457, 12'h557, 12'h557, 12'h457, 12'h557, 12'h457, 12'h447, 12'h447, 12'h446, 12'h346, 12'h346, 12'h346, 12'h447, 12'h447, 12'h457, 12'h557, 12'h557, 12'h557, 12'h457, 12'h457, 12'h457, 12'h457, 12'h557, 12'h557, 12'h557, 
12'h557, 12'h557, 12'h557, 12'h457, 12'h446, 12'h446, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h345, 12'h345, 12'h345, 12'h346, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h556, 12'h567, 12'h678, 12'h779, 12'h889, 12'h89a, 12'h899, 12'h889, 12'h789, 12'h789, 12'h678, 12'h678, 12'h678, 12'h578, 12'h678, 12'h678, 12'h678, 12'h678, 12'h668, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h456, 12'h445, 12'h345, 12'h345, 12'h335, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h334, 12'h334, 12'h334, 12'h234, 12'h234, 12'h344, 12'h344, 12'h334, 12'h334, 12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h334, 12'h233, 12'h233, 12'h222, 12'h122, 12'h112, 
12'h122, 12'h022, 12'h022, 12'h022, 12'h123, 12'h123, 12'h233, 12'h334, 12'h444, 12'h556, 12'h677, 12'h788, 12'h999, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccb, 12'haaa, 12'h988, 12'h766, 12'h555, 12'h444, 12'h444, 12'h344, 12'h334, 12'h334, 12'h345, 12'h456, 12'h566, 12'h667, 12'h677, 12'h778, 12'h789, 12'h99a, 12'haab, 12'haab, 12'h9aa, 12'h89a, 12'h778, 12'h667, 12'h567, 12'h456, 12'h446, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h335, 12'h235, 12'h235, 12'h335, 12'h335, 12'h345, 12'h346, 12'h346, 12'h456, 12'h456, 12'h457, 12'h557, 12'h457, 12'h446, 12'h446, 12'h457, 12'h457, 12'h557, 12'h557, 12'h557, 12'h557, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h557, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h668, 12'h668, 12'h668, 
12'h678, 12'h678, 12'h668, 12'h668, 12'h568, 12'h567, 12'h557, 12'h457, 12'h457, 12'h447, 12'h446, 12'h346, 12'h346, 12'h346, 12'h446, 12'h456, 12'h456, 12'h456, 12'h456, 12'h457, 12'h557, 12'h667, 12'h778, 12'h889, 12'h99a, 12'h99a, 12'h9ab, 12'h9ab, 12'h99a, 12'h89a, 12'h89a, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h678, 12'h678, 12'h668, 12'h668, 12'h678, 12'h678, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h678, 12'h677, 12'h667, 12'h667, 12'h566, 12'h556, 12'h566, 12'h566, 12'h566, 12'h566, 12'h566, 12'h556, 12'h556, 12'h556, 12'h556, 12'h555, 12'h455, 12'h455, 12'h445, 12'h344, 12'h334, 12'h234, 12'h233, 12'h123, 
12'h023, 12'h012, 12'h002, 12'h002, 12'h112, 12'h123, 12'h123, 12'h223, 12'h334, 12'h445, 12'h666, 12'h777, 12'h888, 12'h99a, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heed, 12'hdcc, 12'hbbb, 12'haa9, 12'h887, 12'h666, 12'h555, 12'h444, 12'h344, 12'h344, 12'h334, 12'h234, 12'h345, 12'h556, 12'h567, 12'h677, 12'h678, 12'h678, 12'h778, 12'h99a, 12'habb, 12'haab, 12'h99a, 12'h899, 12'h778, 12'h667, 12'h567, 12'h456, 12'h456, 12'h456, 12'h445, 12'h445, 12'h345, 12'h345, 12'h335, 12'h335, 12'h335, 12'h335, 12'h345, 12'h345, 12'h346, 12'h456, 12'h456, 12'h457, 12'h557, 12'h557, 12'h457, 12'h457, 12'h457, 12'h457, 12'h557, 12'h558, 12'h568, 12'h568, 12'h568, 12'h568, 12'h558, 12'h458, 12'h458, 12'h458, 12'h458, 12'h458, 12'h558, 12'h558, 12'h568, 12'h668, 12'h668, 12'h668, 12'h668, 12'h669, 12'h669, 12'h679, 12'h779, 12'h779, 12'h78a, 
12'h88a, 12'h88a, 12'h88a, 12'h789, 12'h779, 12'h779, 12'h679, 12'h668, 12'h568, 12'h557, 12'h457, 12'h446, 12'h346, 12'h346, 12'h346, 12'h446, 12'h446, 12'h446, 12'h346, 12'h446, 12'h446, 12'h557, 12'h678, 12'h789, 12'h99a, 12'h9ab, 12'habc, 12'habc, 12'haac, 12'h9ab, 12'h99b, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h99b, 12'h9ab, 12'h99b, 12'h89a, 12'h89a, 12'h88a, 12'h789, 12'h789, 12'h889, 12'h89a, 12'h99a, 12'h9aa, 12'h9ab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'h9aa, 12'h99a, 12'h89a, 12'h889, 12'h789, 12'h788, 12'h788, 12'h788, 12'h788, 12'h788, 12'h788, 12'h788, 12'h778, 12'h778, 12'h778, 12'h778, 12'h778, 12'h677, 12'h667, 12'h667, 12'h566, 12'h556, 12'h456, 12'h455, 
12'h345, 12'h334, 12'h234, 12'h334, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h556, 12'h667, 12'h777, 12'h888, 12'h999, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'h999, 12'h777, 12'h555, 12'h444, 12'h333, 12'h333, 12'h334, 12'h223, 12'h223, 12'h334, 12'h456, 12'h567, 12'h678, 12'h678, 12'h678, 12'h778, 12'h99a, 12'habb, 12'habb, 12'h99a, 12'h889, 12'h678, 12'h567, 12'h567, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h335, 12'h335, 12'h335, 12'h345, 12'h346, 12'h446, 12'h456, 12'h457, 12'h557, 12'h567, 12'h567, 12'h557, 12'h457, 12'h457, 12'h557, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h569, 12'h569, 12'h679, 12'h679, 12'h779, 12'h679, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h88a, 12'h88a, 12'h89a, 
12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h89a, 12'h89a, 12'h88a, 12'h88a, 12'h779, 12'h679, 12'h668, 12'h568, 12'h568, 12'h558, 12'h558, 12'h557, 12'h557, 12'h447, 12'h346, 12'h346, 12'h346, 12'h457, 12'h668, 12'h779, 12'h88a, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'habc, 12'h9ab, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ab, 12'h9ab, 12'haac, 12'haac, 12'h9ab, 12'h9ab, 12'h99b, 12'h89a, 12'h89a, 12'h89a, 12'h99a, 12'h9ab, 12'haab, 12'haab, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'habc, 12'habb, 12'haab, 12'h9ab, 12'h89a, 12'h89a, 12'h89a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h899, 12'h889, 12'h889, 12'h788, 
12'h778, 12'h678, 12'h678, 12'h778, 12'h778, 12'h678, 12'h667, 12'h678, 12'h778, 12'h778, 12'h888, 12'h889, 12'h899, 12'h99a, 12'habb, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h998, 12'h776, 12'h544, 12'h433, 12'h333, 12'h333, 12'h334, 12'h223, 12'h113, 12'h334, 12'h456, 12'h567, 12'h667, 12'h668, 12'h678, 12'h778, 12'h99a, 12'haab, 12'haab, 12'h99a, 12'h889, 12'h678, 12'h567, 12'h567, 12'h457, 12'h456, 12'h456, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h346, 12'h346, 12'h456, 12'h457, 12'h557, 12'h567, 12'h568, 12'h568, 12'h557, 12'h558, 12'h568, 12'h568, 12'h568, 12'h669, 12'h669, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h77a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h89b, 12'h99b, 
12'h99b, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h789, 12'h779, 12'h669, 12'h558, 12'h447, 12'h447, 12'h336, 12'h447, 12'h558, 12'h669, 12'h88a, 12'h99b, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'h9ac, 12'h89b, 12'h89a, 12'h79a, 12'h89b, 12'h9ab, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'haac, 12'h9ab, 12'h9ab, 12'h89b, 12'h89b, 12'h9ab, 12'haac, 12'haab, 12'haab, 12'haab, 12'habc, 12'hbbc, 12'hbcd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbcc, 12'hbbc, 12'habc, 12'h9ab, 12'h9ab, 12'haab, 12'haab, 12'haab, 12'hbbb, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hbcc, 12'hbcc, 12'hbcc, 12'hbcc, 12'hbbc, 12'hbbc, 12'habb, 12'haab, 
12'h9aa, 12'h99a, 12'h99a, 12'haab, 12'haab, 12'h99a, 12'h89a, 12'h99a, 12'h99a, 12'h99a, 12'h9aa, 12'h99a, 12'h99a, 12'haab, 12'hbbb, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'ha99, 12'h888, 12'h766, 12'h555, 12'h444, 12'h333, 12'h334, 12'h334, 12'h223, 12'h123, 12'h334, 12'h456, 12'h556, 12'h567, 12'h567, 12'h667, 12'h778, 12'h89a, 12'h9aa, 12'h9aa, 12'h99a, 12'h889, 12'h678, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h346, 12'h346, 12'h345, 12'h345, 12'h346, 12'h346, 12'h346, 12'h457, 12'h557, 12'h568, 12'h668, 12'h568, 12'h568, 12'h568, 12'h568, 12'h668, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h77a, 12'h78a, 12'h78a, 12'h78a, 12'h88a, 12'h78a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 
12'h99c, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'h9ab, 12'h9ab, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h779, 12'h558, 12'h447, 12'h447, 12'h347, 12'h447, 12'h668, 12'h88a, 12'h89a, 12'h89b, 12'h9ac, 12'habc, 12'habc, 12'h9ac, 12'h89b, 12'h78a, 12'h78a, 12'h79a, 12'h9ab, 12'h9bc, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'h9ac, 12'h89b, 12'h89b, 12'h9ab, 12'haac, 12'h9ac, 12'h9ab, 12'h9ab, 12'haac, 12'habc, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcdd, 12'hcdd, 12'hccd, 12'hccd, 12'hccd, 12'hbbc, 12'hbbc, 
12'hbbc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'haab, 12'haab, 12'haab, 12'haab, 12'habc, 12'hbbc, 12'hbbc, 12'habb, 12'hbbb, 12'hbbc, 12'hccc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heed, 12'hdcc, 12'hbba, 12'h998, 12'h887, 12'h766, 12'h655, 12'h544, 12'h444, 12'h334, 12'h334, 12'h223, 12'h224, 12'h335, 12'h456, 12'h556, 12'h456, 12'h557, 12'h667, 12'h778, 12'h889, 12'h99a, 12'h99a, 12'h89a, 12'h889, 12'h678, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h446, 12'h445, 12'h345, 12'h345, 12'h345, 12'h346, 12'h346, 12'h346, 12'h336, 12'h336, 12'h346, 12'h346, 12'h457, 12'h557, 12'h668, 12'h678, 12'h668, 12'h568, 12'h568, 12'h569, 12'h679, 12'h679, 12'h679, 12'h679, 12'h77a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 
12'haac, 12'haac, 12'haac, 12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'h99b, 12'h88a, 12'h88a, 12'h779, 12'h669, 12'h669, 12'h669, 12'h77a, 12'h98b, 12'h99b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h79b, 12'h78a, 12'h78b, 12'h89b, 12'h9ac, 12'habc, 12'habc, 12'habd, 12'habc, 12'habd, 12'habd, 12'habc, 12'h9ab, 12'h99b, 12'h9ab, 12'haac, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'habc, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbcd, 12'hbbc, 12'hbbc, 12'hbbc, 
12'hbbc, 12'hbbc, 12'hbbc, 12'hbcd, 12'hbbc, 12'hbbc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcd, 12'hbcd, 12'hbcc, 12'hbbc, 12'hccc, 12'hccd, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hedd, 12'hccc, 12'hbaa, 12'h888, 12'h877, 12'h766, 12'h555, 12'h444, 12'h333, 12'h334, 12'h334, 12'h223, 12'h223, 12'h335, 12'h446, 12'h556, 12'h456, 12'h557, 12'h667, 12'h678, 12'h889, 12'h89a, 12'h99a, 12'h89a, 12'h789, 12'h678, 12'h567, 12'h557, 12'h557, 12'h456, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h446, 12'h457, 12'h568, 12'h668, 12'h679, 12'h669, 12'h669, 12'h669, 12'h679, 12'h679, 12'h679, 12'h77a, 12'h78a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 
12'haad, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbc, 12'haac, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h88a, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h8ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h78b, 12'h78b, 12'h89b, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habc, 12'habd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'habc, 12'habc, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'habc, 12'habd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 12'hbcd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 
12'hbbc, 12'hbbd, 12'hccd, 12'hccd, 12'hbcd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h887, 12'h776, 12'h666, 12'h554, 12'h444, 12'h333, 12'h333, 12'h334, 12'h223, 12'h224, 12'h335, 12'h446, 12'h556, 12'h456, 12'h557, 12'h567, 12'h678, 12'h789, 12'h889, 12'h89a, 12'h889, 12'h779, 12'h668, 12'h557, 12'h557, 12'h457, 12'h556, 12'h556, 12'h456, 12'h456, 12'h446, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h346, 12'h446, 12'h446, 12'h457, 12'h557, 12'h568, 12'h668, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h77a, 12'h78a, 12'h78a, 12'h78a, 12'h78b, 12'h88b, 12'h89b, 12'h89b, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h89c, 12'h99c, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 
12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbce, 12'hbce, 12'hbbd, 12'hbbd, 12'hbcd, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbc, 12'haac, 12'haac, 12'h99b, 12'h99b, 12'h99b, 12'ha9c, 12'h9ac, 12'h9ac, 12'h8ac, 12'h8ac, 12'h9ac, 12'h9ac, 12'h8ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'habc, 12'habd, 12'habd, 12'habd, 12'habc, 12'haac, 12'h9ac, 12'h9ac, 12'habc, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'habd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbc, 12'hbbc, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 
12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hccb, 12'haa9, 12'h887, 12'h776, 12'h665, 12'h554, 12'h444, 12'h333, 12'h333, 12'h233, 12'h223, 12'h224, 12'h335, 12'h446, 12'h456, 12'h456, 12'h556, 12'h567, 12'h667, 12'h778, 12'h889, 12'h889, 12'h789, 12'h778, 12'h567, 12'h457, 12'h456, 12'h456, 12'h556, 12'h556, 12'h556, 12'h456, 12'h446, 12'h446, 12'h446, 12'h346, 12'h446, 12'h446, 12'h446, 12'h456, 12'h457, 12'h557, 12'h557, 12'h568, 12'h568, 12'h669, 12'h669, 12'h679, 12'h679, 12'h679, 12'h67a, 12'h77a, 12'h78a, 12'h78a, 12'h78b, 12'h88b, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 
12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbac, 12'haac, 12'ha9c, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habc, 12'habc, 12'habd, 12'habd, 12'habd, 12'habc, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habc, 12'habc, 12'habc, 12'habd, 12'hbcd, 12'hcce, 12'hcce, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbc, 12'habc, 12'haac, 12'haac, 12'haac, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 
12'hbbc, 12'habc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hbbd, 12'hbcd, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hcbb, 12'haa9, 12'h887, 12'h766, 12'h665, 12'h544, 12'h443, 12'h333, 12'h333, 12'h233, 12'h223, 12'h224, 12'h335, 12'h446, 12'h456, 12'h456, 12'h556, 12'h557, 12'h567, 12'h678, 12'h779, 12'h789, 12'h778, 12'h678, 12'h557, 12'h456, 12'h456, 12'h446, 12'h456, 12'h556, 12'h556, 12'h456, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h457, 12'h557, 12'h557, 12'h557, 12'h568, 12'h568, 12'h568, 12'h568, 12'h669, 12'h669, 12'h679, 12'h679, 12'h67a, 12'h77a, 12'h77a, 12'h78a, 12'h78b, 12'h88b, 12'h89b, 12'h89c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 
12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'haac, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'habd, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbcd, 12'hbce, 12'hbce, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbc, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'habc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 
12'habc, 12'haac, 12'haac, 12'haac, 12'habc, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hccd, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'heed, 12'hddc, 12'hbbb, 12'h999, 12'h777, 12'h766, 12'h655, 12'h544, 12'h433, 12'h333, 12'h333, 12'h333, 12'h223, 12'h224, 12'h334, 12'h445, 12'h446, 12'h456, 12'h456, 12'h557, 12'h567, 12'h668, 12'h778, 12'h778, 12'h678, 12'h667, 12'h557, 12'h446, 12'h446, 12'h446, 12'h456, 12'h556, 12'h556, 12'h456, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h557, 12'h557, 12'h557, 12'h568, 12'h668, 12'h568, 12'h568, 12'h568, 12'h568, 12'h569, 12'h669, 12'h669, 12'h679, 12'h67a, 12'h67a, 12'h77a, 12'h78a, 12'h78b, 12'h88b, 12'h89b, 12'h89c, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 
12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcbd, 12'hbbd, 12'hbbc, 12'haac, 12'habc, 12'hbbd, 12'hbcd, 12'habd, 12'haac, 12'haac, 12'haad, 12'haac, 12'haac, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'habd, 12'hbcd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbc, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'habc, 12'habc, 12'habc, 12'hbbc, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 
12'haac, 12'haab, 12'h9ab, 12'haab, 12'haac, 12'hbbc, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hccd, 12'hccd, 12'hddd, 12'hdee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hedd, 12'hdcc, 12'hbbb, 12'h999, 12'h776, 12'h665, 12'h555, 12'h544, 12'h433, 12'h333, 12'h333, 12'h334, 12'h224, 12'h224, 12'h334, 12'h445, 12'h445, 12'h446, 12'h456, 12'h556, 12'h557, 12'h667, 12'h678, 12'h678, 12'h667, 12'h567, 12'h456, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h456, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h556, 12'h557, 12'h567, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h568, 12'h568, 12'h568, 12'h569, 12'h669, 12'h669, 12'h679, 12'h67a, 12'h77a, 12'h78a, 12'h78b, 12'h78b, 12'h89b, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 
12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdce, 12'hcce, 12'hccd, 12'hcbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbce, 12'hbbd, 12'habd, 12'habc, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbbd, 12'habd, 12'habd, 12'h9ac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habd, 12'habd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbc, 12'habc, 12'haac, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'haab, 12'haab, 12'haac, 12'haac, 12'haac, 12'haac, 
12'haab, 12'h9ab, 12'h99b, 12'h99b, 12'h9ab, 12'haac, 12'habc, 12'haac, 12'haac, 12'habc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbd, 12'habc, 12'habc, 12'hbbc, 12'hbbc, 12'hccd, 12'hcdd, 12'hdde, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hedd, 12'hccc, 12'hbba, 12'h998, 12'h776, 12'h665, 12'h555, 12'h444, 12'h333, 12'h333, 12'h333, 12'h334, 12'h234, 12'h224, 12'h334, 12'h345, 12'h445, 12'h445, 12'h446, 12'h556, 12'h556, 12'h567, 12'h667, 12'h667, 12'h567, 12'h557, 12'h456, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h556, 12'h557, 12'h667, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h568, 12'h569, 12'h569, 12'h669, 12'h669, 12'h679, 12'h67a, 12'h67a, 12'h78a, 12'h78b, 12'h88b, 12'h89c, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 
12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbcd, 12'hbbd, 12'hbbd, 12'habd, 12'habc, 12'habd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'habd, 12'habc, 12'h9ac, 12'h99c, 12'h99b, 12'h89b, 12'h99b, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'habc, 12'habd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbc, 12'habc, 12'habc, 12'haac, 12'haab, 12'h9ab, 12'h99b, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 
12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ab, 12'haab, 12'haac, 12'habc, 12'hbbc, 12'hbbd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'hbbc, 12'hbbc, 12'hccd, 12'hddd, 12'hdee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h998, 12'h776, 12'h665, 12'h554, 12'h444, 12'h333, 12'h333, 12'h333, 12'h234, 12'h234, 12'h234, 12'h334, 12'h345, 12'h445, 12'h445, 12'h446, 12'h446, 12'h556, 12'h556, 12'h567, 12'h567, 12'h557, 12'h556, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h556, 12'h557, 12'h567, 12'h668, 12'h678, 12'h779, 12'h779, 12'h679, 12'h679, 12'h679, 12'h679, 12'h669, 12'h569, 12'h669, 12'h679, 12'h67a, 12'h67a, 12'h78a, 12'h78b, 12'h88b, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 
12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hcce, 12'hbce, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habc, 12'habd, 12'hbbd, 12'hbcd, 12'hcce, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 12'hccd, 12'hcce, 12'hcce, 12'hbbd, 12'hbbd, 12'haac, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h9ac, 12'habc, 12'hbbd, 12'hbbd, 12'habd, 12'habc, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'habd, 12'habc, 12'habc, 12'haac, 12'haac, 12'h9ab, 12'h99b, 12'h89a, 12'h88a, 12'h78a, 12'h789, 12'h789, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 
12'h89a, 12'h89b, 12'h89a, 12'h88a, 12'h88a, 12'h89a, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'haac, 12'haac, 12'hbbc, 12'hbbc, 12'haac, 12'haab, 12'haab, 12'haab, 12'habc, 12'hbcc, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'haaa, 12'h888, 12'h776, 12'h665, 12'h554, 12'h444, 12'h333, 12'h333, 12'h333, 12'h334, 12'h234, 12'h234, 12'h234, 12'h335, 12'h445, 12'h445, 12'h445, 12'h446, 12'h456, 12'h556, 12'h556, 12'h556, 12'h556, 12'h556, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h446, 12'h557, 12'h567, 12'h668, 12'h678, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h679, 12'h669, 12'h569, 12'h669, 12'h679, 12'h67a, 12'h67a, 12'h78a, 12'h78b, 12'h88b, 12'h89c, 12'h89c, 12'h99c, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 
12'hbce, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hcce, 12'hcde, 12'hcde, 12'hccd, 12'hbbd, 12'habc, 12'h9ac, 12'h99b, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'habd, 12'hbcd, 12'hbcd, 12'habd, 12'h9ac, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'habd, 12'habd, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ab, 12'h99b, 12'h89a, 12'h78a, 12'h789, 12'h679, 12'h679, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h679, 
12'h789, 12'h78a, 12'h78a, 12'h789, 12'h789, 12'h78a, 12'h88a, 12'h88a, 12'h89a, 12'h89a, 12'h99b, 12'h9ab, 12'haab, 12'haac, 12'haab, 12'h9ab, 12'h9ab, 12'h9ab, 12'haab, 12'habc, 12'hbcc, 12'hcdd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccb, 12'haaa, 12'h888, 12'h766, 12'h555, 12'h444, 12'h443, 12'h333, 12'h333, 12'h334, 12'h334, 12'h234, 12'h234, 12'h234, 12'h334, 12'h335, 12'h345, 12'h445, 12'h445, 12'h446, 12'h446, 12'h556, 12'h556, 12'h556, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h335, 12'h335, 12'h435, 12'h446, 12'h456, 12'h557, 12'h667, 12'h668, 12'h779, 12'h779, 12'h789, 12'h78a, 12'h78a, 12'h779, 12'h669, 12'h569, 12'h569, 12'h669, 12'h67a, 12'h67a, 12'h77a, 12'h78b, 12'h88b, 12'h89c, 12'h89c, 12'h99c, 12'h9ad, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hcce, 12'hbcd, 12'hbbd, 12'haac, 12'haac, 12'h99b, 12'h99b, 12'h99b, 12'h9ac, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbbd, 12'h9ac, 12'h88b, 12'h78a, 12'h89b, 12'h99b, 12'h9ac, 12'habc, 12'haac, 12'haac, 12'haab, 12'haac, 12'haab, 12'h9ab, 12'h99b, 12'h89a, 12'h78a, 12'h779, 12'h679, 12'h668, 12'h678, 12'h668, 12'h678, 12'h668, 12'h668, 12'h568, 
12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h779, 12'h789, 12'h78a, 12'h78a, 12'h88a, 12'h89a, 12'h89a, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h9ab, 12'h9ab, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccb, 12'haa9, 12'h888, 12'h666, 12'h555, 12'h444, 12'h343, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h234, 12'h234, 12'h334, 12'h334, 12'h335, 12'h345, 12'h445, 12'h445, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h335, 12'h335, 12'h335, 12'h335, 12'h446, 12'h456, 12'h557, 12'h668, 12'h779, 12'h779, 12'h889, 12'h88a, 12'h88a, 12'h77a, 12'h669, 12'h569, 12'h569, 12'h669, 12'h67a, 12'h67a, 12'h77a, 12'h78b, 12'h88b, 12'h89c, 12'h99c, 12'h99c, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'h99b, 12'h99b, 12'h99b, 12'habc, 12'hbbd, 12'hbcd, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h88b, 12'h89b, 12'h89b, 12'h99b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h89a, 12'h78a, 12'h789, 12'h679, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h468, 
12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h679, 12'h779, 12'h789, 12'h789, 12'h789, 12'h789, 12'h789, 12'h88a, 12'h89a, 12'h89a, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ab, 12'habc, 12'hbcc, 12'hcdd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccb, 12'haa9, 12'h887, 12'h666, 12'h555, 12'h444, 12'h343, 12'h333, 12'h333, 12'h334, 12'h344, 12'h334, 12'h334, 12'h234, 12'h234, 12'h334, 12'h334, 12'h335, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h435, 12'h435, 12'h445, 12'h445, 12'h445, 12'h445, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h446, 12'h557, 12'h667, 12'h668, 12'h779, 12'h789, 12'h88a, 12'h88a, 12'h77a, 12'h669, 12'h569, 12'h569, 12'h669, 12'h66a, 12'h67a, 12'h77b, 12'h78b, 12'h88b, 12'h89c, 12'h99c, 12'h99c, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hcde, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'hedf, 12'hdde, 12'hdde, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hbbd, 12'habc, 12'haac, 12'h99b, 12'h99b, 12'haac, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbbd, 12'haac, 12'h99b, 12'h89b, 12'h88b, 12'h88a, 12'h88a, 12'h89b, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h9ab, 12'h99b, 12'h89a, 12'h88a, 12'h789, 12'h679, 12'h678, 12'h568, 12'h568, 12'h467, 12'h457, 12'h457, 12'h457, 
12'h457, 12'h457, 12'h467, 12'h568, 12'h568, 12'h678, 12'h678, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h679, 12'h789, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h9ab, 12'h9bb, 12'hbbc, 12'hccd, 12'hcdd, 12'hdee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hcbb, 12'h999, 12'h887, 12'h666, 12'h555, 12'h444, 12'h333, 12'h233, 12'h333, 12'h334, 12'h344, 12'h334, 12'h334, 12'h234, 12'h234, 12'h234, 12'h334, 12'h335, 12'h435, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h435, 12'h335, 12'h435, 12'h435, 12'h445, 12'h445, 12'h445, 12'h435, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h446, 12'h557, 12'h668, 12'h678, 12'h779, 12'h78a, 12'h78a, 12'h779, 12'h669, 12'h569, 12'h569, 12'h669, 12'h66a, 12'h67a, 12'h77b, 12'h78b, 12'h88b, 12'h89c, 12'h99c, 12'h99d, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haae, 12'habe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'hedf, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'habc, 12'haac, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89a, 12'h89a, 12'h78a, 12'h789, 12'h678, 12'h568, 12'h567, 12'h457, 12'h357, 12'h457, 12'h457, 
12'h457, 12'h457, 12'h457, 12'h467, 12'h568, 12'h568, 12'h568, 12'h568, 12'h678, 12'h678, 12'h568, 12'h678, 12'h678, 12'h789, 12'h88a, 12'h89a, 12'h89a, 12'h88a, 12'h89a, 12'h89a, 12'h9ab, 12'habc, 12'hbcc, 12'hcdd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h887, 12'h666, 12'h555, 12'h444, 12'h333, 12'h233, 12'h233, 12'h334, 12'h344, 12'h344, 12'h334, 12'h234, 12'h224, 12'h224, 12'h334, 12'h334, 12'h335, 12'h445, 12'h335, 12'h335, 12'h435, 12'h435, 12'h445, 12'h445, 12'h435, 12'h435, 12'h334, 12'h334, 12'h334, 12'h435, 12'h445, 12'h445, 12'h435, 12'h435, 12'h335, 12'h335, 12'h335, 12'h335, 12'h346, 12'h447, 12'h557, 12'h668, 12'h668, 12'h779, 12'h779, 12'h679, 12'h669, 12'h669, 12'h669, 12'h669, 12'h67a, 12'h67a, 12'h78b, 12'h78b, 12'h89c, 12'h89c, 12'h99c, 12'h9ad, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'habe, 12'habe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'heef, 12'heef, 12'hede, 12'hede, 12'hdde, 12'hede, 12'hedf, 12'heef, 12'heef, 12'hedf, 12'hddf, 12'hedf, 12'hddf, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h789, 12'h679, 12'h568, 12'h467, 12'h457, 12'h357, 12'h357, 12'h357, 
12'h357, 12'h357, 12'h357, 12'h457, 12'h457, 12'h457, 12'h457, 12'h467, 12'h568, 12'h568, 12'h568, 12'h568, 12'h568, 12'h679, 12'h789, 12'h89a, 12'h789, 12'h789, 12'h78a, 12'h89a, 12'h9ab, 12'habb, 12'hbcc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h887, 12'h666, 12'h554, 12'h343, 12'h233, 12'h223, 12'h233, 12'h334, 12'h344, 12'h344, 12'h334, 12'h334, 12'h224, 12'h224, 12'h224, 12'h334, 12'h335, 12'h435, 12'h335, 12'h335, 12'h335, 12'h435, 12'h435, 12'h445, 12'h435, 12'h334, 12'h324, 12'h324, 12'h324, 12'h334, 12'h435, 12'h445, 12'h445, 12'h445, 12'h335, 12'h335, 12'h325, 12'h225, 12'h335, 12'h446, 12'h447, 12'h557, 12'h568, 12'h668, 12'h669, 12'h669, 12'h669, 12'h669, 12'h669, 12'h66a, 12'h67a, 12'h67a, 12'h78b, 12'h88b, 12'h89c, 12'h89c, 12'h99c, 12'h9ad, 12'h9ad, 12'haad, 12'haad, 12'habe, 12'habe, 12'habe, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hbce, 12'hcce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hedf, 12'heef, 12'heef, 12'heef, 12'hede, 12'hede, 12'hede, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'haac, 12'habd, 12'hbbd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h99b, 12'h89b, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h89a, 12'h88a, 12'h78a, 12'h779, 12'h678, 12'h568, 12'h457, 12'h457, 12'h457, 12'h457, 
12'h457, 12'h457, 12'h457, 12'h457, 12'h457, 12'h446, 12'h346, 12'h456, 12'h457, 12'h557, 12'h567, 12'h567, 12'h667, 12'h678, 12'h788, 12'h789, 12'h789, 12'h789, 12'h789, 12'h89a, 12'h99a, 12'haab, 12'hbbc, 12'hbcc, 12'hcdd, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h777, 12'h666, 12'h554, 12'h443, 12'h233, 12'h222, 12'h223, 12'h334, 12'h344, 12'h344, 12'h334, 12'h334, 12'h234, 12'h224, 12'h224, 12'h334, 12'h335, 12'h335, 12'h334, 12'h334, 12'h334, 12'h334, 12'h434, 12'h434, 12'h434, 12'h334, 12'h324, 12'h323, 12'h324, 12'h334, 12'h434, 12'h435, 12'h445, 12'h445, 12'h335, 12'h335, 12'h325, 12'h225, 12'h335, 12'h336, 12'h446, 12'h457, 12'h557, 12'h568, 12'h568, 12'h669, 12'h669, 12'h679, 12'h679, 12'h67a, 12'h67a, 12'h77a, 12'h78b, 12'h88b, 12'h89c, 12'h99c, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habe, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hbbd, 12'hbbc, 12'habc, 12'habd, 12'habd, 12'hbbd, 12'habd, 12'haad, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ab, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h78a, 12'h779, 12'h679, 12'h669, 12'h668, 12'h558, 12'h557, 12'h557, 
12'h557, 12'h557, 12'h557, 12'h556, 12'h556, 12'h446, 12'h445, 12'h445, 12'h446, 12'h556, 12'h556, 12'h566, 12'h667, 12'h667, 12'h778, 12'h778, 12'h778, 12'h778, 12'h889, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hbcc, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hbbb, 12'h999, 12'h877, 12'h666, 12'h554, 12'h443, 12'h333, 12'h322, 12'h333, 12'h333, 12'h444, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h434, 12'h434, 12'h333, 12'h333, 12'h333, 12'h333, 12'h434, 12'h434, 12'h434, 12'h434, 12'h334, 12'h334, 12'h334, 12'h335, 12'h235, 12'h335, 12'h336, 12'h346, 12'h447, 12'h557, 12'h568, 12'h668, 12'h669, 12'h679, 12'h679, 12'h67a, 12'h67a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 
12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'haad, 12'h9ad, 12'h9ac, 12'h9ac, 12'h9ac, 12'h9ac, 12'h89b, 12'h88b, 12'h78a, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h779, 12'h779, 12'h679, 12'h669, 12'h668, 12'h558, 12'h557, 12'h557, 
12'h557, 12'h557, 12'h557, 12'h556, 12'h546, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h556, 12'h666, 12'h667, 12'h667, 12'h677, 12'h777, 12'h778, 12'h778, 12'h889, 12'h99a, 12'h9ab, 12'habb, 12'hbbc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hbbb, 12'h998, 12'h877, 12'h666, 12'h554, 12'h444, 12'h333, 12'h322, 12'h333, 12'h433, 12'h434, 12'h334, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h434, 12'h434, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h234, 12'h235, 12'h335, 12'h346, 12'h447, 12'h457, 12'h568, 12'h668, 12'h679, 12'h679, 12'h77a, 12'h77a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h89c, 12'h9ac, 12'h9ac, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 
12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hcde, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'habd, 12'haad, 12'h9ad, 12'h99c, 12'h99c, 12'h9ac, 12'h89c, 12'h89b, 12'h89b, 12'h78b, 12'h78a, 12'h77a, 12'h67a, 12'h679, 12'h669, 12'h669, 12'h668, 12'h568, 12'h558, 12'h557, 12'h557, 12'h547, 
12'h547, 12'h557, 12'h556, 12'h546, 12'h546, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h556, 12'h566, 12'h666, 12'h666, 12'h667, 12'h777, 12'h778, 12'h789, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccc, 12'hcdd, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hbbb, 12'h998, 12'h877, 12'h665, 12'h544, 12'h443, 12'h433, 12'h322, 12'h322, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h234, 12'h235, 12'h335, 12'h346, 12'h447, 12'h557, 12'h568, 12'h668, 12'h679, 12'h679, 12'h77a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h89b, 12'h9ac, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 
12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hbce, 12'hbbd, 12'habd, 12'haad, 12'h99c, 12'h99c, 12'h89c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h78b, 12'h78a, 12'h679, 12'h569, 12'h568, 12'h558, 12'h558, 12'h558, 12'h557, 12'h557, 12'h447, 12'h446, 
12'h446, 12'h546, 12'h546, 12'h546, 12'h546, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h555, 12'h556, 12'h566, 12'h666, 12'h667, 12'h778, 12'h778, 12'h889, 12'h99a, 12'haab, 12'hbbb, 12'hbcc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hbba, 12'h988, 12'h777, 12'h665, 12'h544, 12'h443, 12'h433, 12'h322, 12'h322, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h234, 12'h235, 12'h335, 12'h346, 12'h447, 12'h557, 12'h568, 12'h668, 12'h679, 12'h77a, 12'h78a, 12'h78a, 12'h88b, 12'h89b, 12'h99c, 12'h9ac, 12'h9ac, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 
12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hede, 12'hede, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hbce, 12'hbbd, 12'haad, 12'haac, 12'h99c, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78a, 12'h679, 12'h569, 12'h558, 12'h458, 12'h458, 12'h457, 12'h557, 12'h557, 12'h447, 12'h446, 
12'h446, 12'h446, 12'h446, 12'h446, 12'h546, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h435, 12'h445, 12'h445, 12'h445, 12'h445, 12'h556, 12'h556, 12'h666, 12'h677, 12'h778, 12'h889, 12'h99a, 12'h9ab, 12'habb, 12'hbcc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heee, 12'hddc, 12'hbba, 12'h988, 12'h776, 12'h665, 12'h554, 12'h443, 12'h433, 12'h322, 12'h322, 12'h322, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h324, 12'h324, 12'h224, 12'h224, 12'h235, 12'h335, 12'h336, 12'h447, 12'h457, 12'h568, 12'h668, 12'h679, 12'h78a, 12'h88a, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hcbd, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hdde, 12'hcde, 12'hcce, 12'hbbd, 12'hbbd, 12'haac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78a, 12'h679, 12'h669, 12'h558, 12'h458, 12'h458, 12'h457, 12'h457, 12'h457, 12'h447, 12'h446, 
12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h546, 12'h546, 12'h445, 12'h445, 12'h435, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h445, 12'h555, 12'h556, 12'h667, 12'h778, 12'h889, 12'h89a, 12'h9aa, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'hddd, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heed, 12'hddc, 12'hbaa, 12'h888, 12'h776, 12'h665, 12'h554, 12'h544, 12'h433, 12'h333, 12'h322, 12'h322, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h323, 12'h324, 12'h324, 12'h224, 12'h224, 12'h225, 12'h335, 12'h336, 12'h447, 12'h457, 12'h568, 12'h668, 12'h679, 12'h78a, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hcde, 12'hcce, 12'hccd, 12'hbbd, 12'haac, 12'h9ac, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h78a, 12'h77a, 12'h679, 12'h669, 12'h568, 12'h558, 12'h558, 12'h557, 12'h557, 12'h557, 12'h547, 
12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h334, 12'h334, 12'h334, 12'h334, 12'h344, 12'h445, 12'h455, 12'h556, 12'h667, 12'h778, 12'h789, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heed, 12'hddc, 12'hbaa, 12'h888, 12'h766, 12'h665, 12'h544, 12'h544, 12'h433, 12'h333, 12'h322, 12'h322, 12'h322, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h323, 12'h323, 12'h324, 12'h224, 12'h224, 12'h225, 12'h335, 12'h336, 12'h446, 12'h457, 12'h568, 12'h668, 12'h679, 12'h88a, 12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'haac, 12'haac, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hbbd, 12'haac, 12'h9ac, 12'h99c, 12'h89b, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h77a, 12'h679, 12'h669, 12'h668, 12'h558, 12'h558, 12'h557, 12'h557, 12'h557, 
12'h547, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h435, 12'h334, 12'h334, 12'h334, 12'h334, 12'h445, 12'h445, 12'h555, 12'h556, 12'h667, 12'h778, 12'h789, 12'h89a, 12'h9aa, 12'habb, 12'hbcc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heed, 12'hddc, 12'hbaa, 12'h887, 12'h766, 12'h655, 12'h544, 12'h443, 12'h433, 12'h332, 12'h322, 12'h322, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h224, 12'h224, 12'h224, 12'h224, 12'h235, 12'h336, 12'h446, 12'h457, 12'h568, 12'h668, 12'h679, 12'h88a, 12'h89b, 12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 
12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hdde, 12'hcde, 12'hcce, 12'hbbd, 12'haac, 12'h9ac, 12'h99b, 12'h89b, 12'h78a, 12'h78a, 12'h78a, 12'h77a, 12'h779, 12'h679, 12'h668, 12'h568, 12'h558, 12'h557, 12'h557, 12'h557, 
12'h557, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h435, 12'h334, 12'h334, 12'h334, 12'h334, 12'h345, 12'h445, 12'h445, 12'h456, 12'h567, 12'h668, 12'h778, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heed, 12'hddc, 12'hbaa, 12'h887, 12'h766, 12'h655, 12'h544, 12'h444, 12'h433, 12'h333, 12'h333, 12'h323, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h433, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h224, 12'h224, 12'h224, 12'h224, 12'h235, 12'h336, 12'h446, 12'h457, 12'h558, 12'h668, 12'h679, 12'h78a, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'haac, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 
12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'hfef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hcde, 12'hbce, 12'habd, 12'haac, 12'h9ac, 12'h89b, 12'h88b, 12'h78a, 12'h78a, 12'h77a, 12'h779, 12'h669, 12'h668, 12'h558, 12'h558, 12'h557, 12'h557, 12'h557, 
12'h557, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h435, 12'h335, 12'h334, 12'h334, 12'h344, 12'h345, 12'h445, 12'h445, 12'h445, 12'h456, 12'h567, 12'h778, 12'h889, 12'h89a, 12'haab, 12'hbbc, 12'hccc, 12'hcdd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heed, 12'hddc, 12'hbaa, 12'h887, 12'h766, 12'h554, 12'h544, 12'h443, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h224, 12'h224, 12'h224, 12'h224, 12'h225, 12'h336, 12'h346, 12'h457, 12'h558, 12'h568, 12'h679, 12'h78a, 12'h88a, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h89b, 12'h88b, 12'h89b, 12'h89b, 12'h89c, 12'h99c, 12'h99c, 12'haac, 12'haad, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 
12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hcde, 12'hbce, 12'hbbd, 12'habd, 12'h9ac, 12'h99b, 12'h88b, 12'h78a, 12'h77a, 12'h779, 12'h669, 12'h668, 12'h568, 12'h558, 12'h557, 12'h557, 12'h557, 
12'h547, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h446, 12'h567, 12'h678, 12'h789, 12'h89a, 12'h9aa, 12'hbbb, 12'hbcc, 12'hcdd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfee, 12'heed, 12'hdcc, 12'hbaa, 12'h887, 12'h666, 12'h554, 12'h543, 12'h443, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h224, 12'h224, 12'h224, 12'h224, 12'h225, 12'h235, 12'h346, 12'h457, 12'h558, 12'h568, 12'h669, 12'h779, 12'h78a, 12'h78a, 12'h78a, 12'h88b, 12'h88b, 12'h88b, 12'h78b, 12'h88b, 12'h88b, 12'h88b, 12'h89c, 12'h99c, 12'h99c, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hcce, 12'hcce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hcde, 12'hcce, 12'hbcd, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h78a, 12'h779, 12'h669, 12'h668, 12'h568, 12'h558, 12'h557, 12'h557, 12'h557, 
12'h447, 12'h446, 12'h446, 12'h446, 12'h446, 12'h436, 12'h435, 12'h335, 12'h335, 12'h435, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h345, 12'h345, 12'h556, 12'h678, 12'h889, 12'h89a, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfee, 12'heed, 12'hddc, 12'hbaa, 12'h887, 12'h666, 12'h544, 12'h443, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h224, 12'h224, 12'h224, 12'h224, 12'h225, 12'h235, 12'h336, 12'h447, 12'h557, 12'h558, 12'h669, 12'h679, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h78b, 12'h88b, 12'h88b, 12'h99c, 12'h99c, 12'h99c, 12'h9ac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hcde, 12'hcce, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h779, 12'h679, 12'h669, 12'h668, 12'h568, 12'h558, 12'h557, 12'h457, 
12'h447, 12'h446, 12'h446, 12'h446, 12'h446, 12'h436, 12'h335, 12'h335, 12'h335, 12'h435, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h345, 12'h344, 12'h344, 12'h335, 12'h335, 12'h456, 12'h668, 12'h789, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfee, 12'heed, 12'hddc, 12'hbaa, 12'h887, 12'h766, 12'h544, 12'h433, 12'h433, 12'h433, 12'h333, 12'h433, 12'h433, 12'h434, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h323, 12'h224, 12'h224, 12'h224, 12'h224, 12'h225, 12'h235, 12'h336, 12'h447, 12'h457, 12'h558, 12'h568, 12'h669, 12'h679, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h78b, 12'h88b, 12'h88b, 12'h89c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'habd, 12'hbbd, 
12'hbcd, 12'hbcd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hdde, 12'hcce, 12'hbbd, 12'haac, 12'h9ab, 12'h89a, 12'h88a, 12'h789, 12'h779, 12'h669, 12'h668, 12'h558, 12'h557, 
12'h557, 12'h447, 12'h446, 12'h446, 12'h446, 12'h446, 12'h335, 12'h335, 12'h335, 12'h335, 12'h345, 12'h345, 12'h345, 12'h445, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h335, 12'h446, 12'h667, 12'h778, 12'h789, 12'h89a, 12'h9aa, 12'habb, 12'hbcc, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heed, 12'hdcc, 12'hbaa, 12'h877, 12'h765, 12'h544, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h324, 12'h224, 12'h224, 12'h224, 12'h225, 12'h225, 12'h336, 12'h446, 12'h457, 12'h558, 12'h568, 12'h669, 12'h679, 12'h77a, 12'h78a, 12'h88a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h88b, 12'h78b, 12'h78a, 12'h78b, 12'h88b, 12'h88b, 12'h89b, 12'h99c, 12'haac, 12'haac, 
12'habd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hedf, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hcce, 12'hbcd, 12'hbbc, 12'haac, 12'h99b, 12'h89a, 12'h88a, 12'h779, 12'h679, 12'h668, 12'h558, 
12'h557, 12'h447, 12'h447, 12'h446, 12'h446, 12'h446, 12'h346, 12'h435, 12'h335, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h335, 12'h345, 12'h556, 12'h667, 12'h778, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'heed, 12'hdcc, 12'haaa, 12'h877, 12'h665, 12'h544, 12'h433, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h323, 12'h334, 12'h324, 12'h224, 12'h224, 12'h225, 12'h225, 12'h336, 12'h446, 12'h447, 12'h558, 12'h568, 12'h669, 12'h779, 12'h77a, 12'h88a, 12'h88b, 12'h89b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h88b, 12'h77b, 12'h77a, 12'h67a, 12'h67a, 12'h77a, 12'h77a, 12'h78a, 12'h88b, 12'h99b, 12'h9ac, 
12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbcd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hcde, 12'hccd, 12'hbbd, 12'haac, 12'haab, 12'h99b, 12'h88a, 12'h779, 12'h679, 12'h668, 
12'h557, 12'h557, 12'h447, 12'h447, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h556, 12'h667, 12'h678, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hedd, 12'hdcc, 12'haaa, 12'h877, 12'h655, 12'h544, 12'h443, 12'h443, 12'h433, 12'h433, 12'h433, 12'h333, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h233, 12'h233, 12'h333, 12'h333, 12'h233, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h333, 12'h333, 12'h333, 12'h334, 12'h324, 12'h224, 12'h224, 12'h224, 12'h225, 12'h335, 12'h346, 12'h447, 12'h457, 12'h558, 12'h669, 12'h779, 12'h78a, 12'h88b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h89b, 12'h88b, 12'h88b, 12'h77a, 12'h66a, 12'h569, 12'h569, 12'h569, 12'h569, 12'h679, 12'h78a, 12'h88b, 12'h89b, 
12'h9ac, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hbcd, 12'hbbc, 12'haab, 12'h99a, 12'h88a, 12'h779, 12'h669, 
12'h668, 12'h557, 12'h447, 12'h447, 12'h447, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h446, 12'h556, 12'h667, 12'h788, 12'h99a, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hedd, 12'hccc, 12'haaa, 12'h877, 12'h655, 12'h544, 12'h433, 12'h443, 12'h443, 12'h433, 12'h333, 12'h333, 12'h322, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h333, 12'h333, 12'h333, 12'h334, 12'h324, 12'h224, 12'h224, 12'h224, 12'h225, 12'h235, 12'h346, 12'h447, 12'h457, 12'h558, 12'h669, 12'h77a, 12'h88a, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h99c, 12'h99c, 12'h99c, 12'h99b, 12'h98b, 12'h88b, 12'h88b, 12'h77b, 12'h77a, 12'h669, 12'h569, 12'h559, 12'h559, 12'h459, 12'h569, 12'h679, 12'h77a, 12'h88a, 
12'h89b, 12'h9ab, 12'haac, 12'habc, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hdde, 12'hcce, 12'hccd, 12'hbbc, 12'h9ab, 12'h88a, 12'h88a, 12'h779, 
12'h668, 12'h557, 12'h447, 12'h457, 12'h457, 12'h457, 12'h446, 12'h446, 12'h446, 12'h446, 12'h345, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h345, 12'h445, 12'h446, 12'h556, 12'h667, 12'h778, 12'h899, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hedd, 12'hccc, 12'haa9, 12'h776, 12'h655, 12'h544, 12'h443, 12'h444, 12'h444, 12'h433, 12'h433, 12'h323, 12'h222, 12'h222, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h333, 12'h333, 12'h334, 12'h334, 12'h224, 12'h224, 12'h224, 12'h225, 12'h235, 12'h346, 12'h447, 12'h557, 12'h568, 12'h669, 12'h77a, 12'h88a, 12'h99b, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'h99c, 12'h99c, 12'h99b, 12'h98b, 12'h88b, 12'h88b, 12'h77a, 12'h66a, 12'h569, 12'h459, 12'h458, 12'h458, 12'h458, 12'h569, 12'h679, 12'h67a, 
12'h78a, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hccd, 12'hbbc, 12'h99b, 12'h88a, 12'h779, 
12'h568, 12'h457, 12'h447, 12'h457, 12'h557, 12'h457, 12'h456, 12'h457, 12'h557, 12'h456, 12'h335, 12'h335, 12'h345, 12'h446, 12'h456, 12'h456, 12'h445, 12'h345, 12'h345, 12'h335, 12'h445, 12'h556, 12'h557, 12'h667, 12'h778, 12'h889, 12'h99a, 12'habb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'heee, 12'hedd, 12'hccc, 12'haa9, 12'h776, 12'h655, 12'h544, 12'h544, 12'h444, 12'h444, 12'h444, 12'h433, 12'h323, 12'h212, 12'h222, 12'h223, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h222, 12'h222, 12'h222, 12'h323, 12'h333, 12'h444, 12'h433, 12'h333, 12'h333, 12'h433, 12'h433, 12'h333, 12'h323, 12'h323, 12'h333, 12'h333, 12'h334, 12'h324, 12'h224, 12'h224, 12'h224, 12'h224, 12'h235, 12'h446, 12'h457, 12'h558, 12'h668, 12'h679, 12'h78a, 12'h88b, 12'h99b, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'haad, 12'haad, 12'haac, 12'haac, 12'haac, 12'h99c, 12'h99c, 12'h99b, 12'h99b, 12'h88b, 12'h77a, 12'h67a, 12'h569, 12'h559, 12'h458, 12'h348, 12'h348, 12'h458, 12'h558, 12'h569, 
12'h679, 12'h78a, 12'h89b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'heee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hccd, 12'hbbc, 12'haab, 12'h88a, 
12'h779, 12'h668, 12'h558, 12'h557, 12'h557, 12'h557, 12'h567, 12'h567, 12'h557, 12'h456, 12'h346, 12'h335, 12'h346, 12'h446, 12'h456, 12'h456, 12'h445, 12'h345, 12'h345, 12'h334, 12'h335, 12'h556, 12'h556, 12'h667, 12'h778, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hffe, 12'heee, 12'hedd, 12'hdcc, 12'haa9, 12'h776, 12'h665, 12'h655, 12'h554, 12'h544, 12'h443, 12'h444, 12'h444, 12'h333, 12'h212, 12'h222, 12'h223, 12'h233, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h222, 12'h212, 12'h212, 12'h223, 12'h433, 12'h444, 12'h444, 12'h333, 12'h333, 12'h433, 12'h433, 12'h323, 12'h322, 12'h323, 12'h333, 12'h333, 12'h334, 12'h324, 12'h324, 12'h224, 12'h214, 12'h224, 12'h335, 12'h446, 12'h557, 12'h568, 12'h668, 12'h779, 12'h88a, 12'h99b, 12'h99b, 12'haac, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'h99c, 12'h99b, 12'h88b, 12'h77a, 12'h669, 12'h559, 12'h458, 12'h348, 12'h348, 12'h458, 12'h458, 12'h458, 
12'h569, 12'h679, 12'h78a, 12'h88a, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hcde, 12'hccd, 12'hbbd, 12'haac, 
12'h99b, 12'h88a, 12'h779, 12'h668, 12'h668, 12'h668, 12'h779, 12'h678, 12'h667, 12'h557, 12'h446, 12'h346, 12'h446, 12'h456, 12'h446, 12'h445, 12'h345, 12'h345, 12'h345, 12'h334, 12'h334, 12'h445, 12'h556, 12'h667, 12'h667, 12'h788, 12'h999, 12'haaa, 12'hbbc, 12'hccd, 12'hddd, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfee, 12'heee, 12'hedd, 12'hccc, 12'haa9, 12'h776, 12'h665, 12'h654, 12'h544, 12'h433, 12'h433, 12'h444, 12'h444, 12'h333, 12'h222, 12'h222, 12'h223, 12'h233, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h222, 12'h222, 12'h222, 12'h323, 12'h433, 12'h444, 12'h433, 12'h333, 12'h333, 12'h433, 12'h333, 12'h322, 12'h322, 12'h322, 12'h322, 12'h323, 12'h334, 12'h324, 12'h324, 12'h224, 12'h224, 12'h224, 12'h335, 12'h446, 12'h457, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'h99b, 12'h88b, 12'h77a, 12'h669, 12'h558, 12'h348, 12'h348, 12'h458, 12'h458, 12'h458, 
12'h458, 12'h568, 12'h569, 12'h679, 12'h78a, 12'h89b, 12'h9ab, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 
12'hbbc, 12'h9ab, 12'h88a, 12'h779, 12'h668, 12'h779, 12'h88a, 12'h789, 12'h668, 12'h567, 12'h557, 12'h456, 12'h456, 12'h456, 12'h446, 12'h345, 12'h345, 12'h345, 12'h345, 12'h334, 12'h334, 12'h445, 12'h556, 12'h667, 12'h667, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfee, 12'heee, 12'hddd, 12'hccc, 12'ha99, 12'h766, 12'h655, 12'h544, 12'h433, 12'h433, 12'h433, 12'h443, 12'h444, 12'h433, 12'h323, 12'h223, 12'h223, 12'h233, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h223, 12'h222, 12'h223, 12'h333, 12'h433, 12'h444, 12'h333, 12'h333, 12'h322, 12'h332, 12'h322, 12'h322, 12'h322, 12'h222, 12'h222, 12'h323, 12'h324, 12'h334, 12'h324, 12'h224, 12'h224, 12'h224, 12'h335, 12'h346, 12'h457, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h89a, 12'h99b, 12'haac, 12'haac, 12'haac, 12'hbbc, 12'hbbd, 12'hcbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'h99b, 12'h88a, 12'h679, 12'h569, 12'h458, 12'h448, 12'h458, 12'h458, 12'h458, 
12'h357, 12'h347, 12'h347, 12'h558, 12'h679, 12'h78a, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 
12'hccd, 12'hbbc, 12'haab, 12'h78a, 12'h679, 12'h889, 12'h99a, 12'h88a, 12'h778, 12'h668, 12'h567, 12'h557, 12'h557, 12'h557, 12'h456, 12'h345, 12'h345, 12'h345, 12'h345, 12'h334, 12'h445, 12'h445, 12'h556, 12'h667, 12'h677, 12'h778, 12'h889, 12'h9aa, 12'hbbb, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'heee, 12'heed, 12'hddd, 12'hccc, 12'haa9, 12'h776, 12'h655, 12'h543, 12'h432, 12'h433, 12'h433, 12'h443, 12'h444, 12'h433, 12'h333, 12'h333, 12'h333, 12'h233, 12'h233, 12'h233, 12'h233, 12'h233, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h333, 12'h333, 12'h333, 12'h433, 12'h333, 12'h322, 12'h322, 12'h333, 12'h333, 12'h322, 12'h322, 12'h322, 12'h322, 12'h323, 12'h334, 12'h334, 12'h334, 12'h324, 12'h324, 12'h225, 12'h335, 12'h346, 12'h446, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h88a, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'hbbc, 12'hbbd, 12'hccd, 12'hccd, 12'hcce, 12'hccd, 12'hcbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'h88b, 12'h77a, 12'h669, 12'h458, 12'h447, 12'h347, 12'h337, 
12'h236, 12'h236, 12'h237, 12'h457, 12'h568, 12'h679, 12'h78a, 12'h88a, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hcde, 12'hccd, 12'hbbc, 12'h89a, 12'h779, 12'h88a, 12'h9ab, 12'h99a, 12'h789, 12'h678, 12'h678, 12'h667, 12'h567, 12'h567, 12'h456, 12'h346, 12'h345, 12'h345, 12'h345, 12'h445, 12'h445, 12'h545, 12'h556, 12'h666, 12'h667, 12'h778, 12'h889, 12'h9aa, 12'hbbb, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'heee, 12'heed, 12'hddd, 12'hccc, 12'haaa, 12'h887, 12'h765, 12'h543, 12'h432, 12'h433, 12'h433, 12'h433, 12'h444, 12'h444, 12'h433, 12'h333, 12'h333, 12'h333, 12'h233, 12'h233, 12'h233, 12'h233, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h322, 12'h333, 12'h433, 12'h433, 12'h433, 12'h323, 12'h323, 12'h323, 12'h333, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h335, 12'h346, 12'h446, 12'h457, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h88a, 12'h99b, 12'h99b, 12'h99b, 12'haab, 12'haac, 12'haac, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hcbd, 12'hbbd, 12'hbbd, 12'haac, 12'h99b, 12'h77a, 12'h668, 12'h458, 12'h337, 12'h236, 
12'h226, 12'h126, 12'h126, 12'h337, 12'h457, 12'h568, 12'h669, 12'h779, 12'h88a, 12'h99b, 12'h99c, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdef, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hcde, 12'hccd, 12'h99b, 12'h78a, 12'h99a, 12'haab, 12'h9ab, 12'h88a, 12'h789, 12'h778, 12'h678, 12'h668, 12'h567, 12'h557, 12'h456, 12'h346, 12'h446, 12'h445, 12'h445, 12'h445, 12'h445, 12'h545, 12'h556, 12'h667, 12'h778, 12'h889, 12'h99a, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 
12'heee, 12'hedd, 12'hddd, 12'hccc, 12'hbaa, 12'h988, 12'h776, 12'h543, 12'h422, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h434, 12'h334, 12'h333, 12'h333, 12'h233, 12'h233, 12'h233, 12'h233, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h433, 12'h444, 12'h444, 12'h434, 12'h434, 12'h433, 12'h333, 12'h334, 12'h434, 12'h434, 12'h435, 12'h335, 12'h335, 12'h335, 12'h335, 12'h336, 12'h446, 12'h446, 12'h557, 12'h568, 12'h668, 12'h779, 12'h789, 12'h88a, 12'h88a, 12'h88a, 12'h99a, 12'h99b, 12'h99b, 12'ha9b, 12'haab, 12'haac, 12'haac, 12'haac, 12'haac, 12'hbac, 12'hbbc, 12'hbbc, 12'hbbc, 12'haac, 12'haac, 12'h99b, 12'h88a, 12'h779, 12'h668, 12'h457, 12'h346, 
12'h236, 12'h236, 12'h126, 12'h236, 12'h347, 12'h457, 12'h558, 12'h669, 12'h779, 12'h88a, 12'h99b, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hcce, 12'haab, 12'h88a, 12'h99a, 12'haab, 12'h9ab, 12'h89a, 12'h88a, 12'h789, 12'h779, 12'h678, 12'h667, 12'h567, 12'h456, 12'h456, 12'h456, 12'h445, 12'h445, 12'h444, 12'h445, 12'h445, 12'h556, 12'h667, 12'h778, 12'h889, 12'h99a, 12'hbbb, 12'hccc, 12'hcdd, 12'hddd, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 
12'heee, 12'hedd, 12'hddd, 12'hccc, 12'hbba, 12'ha99, 12'h877, 12'h554, 12'h432, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h444, 12'h444, 12'h344, 12'h333, 12'h233, 12'h233, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h322, 12'h333, 12'h444, 12'h544, 12'h555, 12'h545, 12'h544, 12'h444, 12'h434, 12'h434, 12'h434, 12'h434, 12'h445, 12'h445, 12'h435, 12'h435, 12'h335, 12'h335, 12'h435, 12'h446, 12'h446, 12'h457, 12'h557, 12'h557, 12'h668, 12'h679, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h98a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'haab, 12'h99b, 12'h99b, 12'h88a, 12'h779, 12'h668, 12'h557, 
12'h447, 12'h346, 12'h236, 12'h236, 12'h347, 12'h347, 12'h457, 12'h558, 12'h669, 12'h779, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'habd, 12'haad, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdef, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hcce, 12'haac, 12'h89a, 12'h99a, 12'h99b, 12'h9ab, 12'h99b, 12'h99a, 12'h889, 12'h789, 12'h678, 12'h668, 12'h567, 12'h556, 12'h456, 12'h456, 12'h456, 12'h445, 12'h445, 12'h444, 12'h445, 12'h556, 12'h667, 12'h778, 12'h889, 12'h999, 12'haab, 12'hbcc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 
12'heee, 12'hedd, 12'hddd, 12'hdcc, 12'hcbb, 12'haa9, 12'h988, 12'h655, 12'h433, 12'h443, 12'h433, 12'h433, 12'h333, 12'h433, 12'h434, 12'h444, 12'h444, 12'h344, 12'h333, 12'h233, 12'h233, 12'h334, 12'h334, 12'h333, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h323, 12'h444, 12'h555, 12'h655, 12'h655, 12'h655, 12'h555, 12'h544, 12'h544, 12'h444, 12'h434, 12'h434, 12'h435, 12'h435, 12'h435, 12'h335, 12'h335, 12'h335, 12'h335, 12'h436, 12'h446, 12'h446, 12'h446, 12'h447, 12'h557, 12'h568, 12'h668, 12'h668, 12'h668, 12'h668, 12'h779, 12'h779, 12'h889, 12'h889, 12'h88a, 12'h88a, 12'h88a, 12'h98a, 12'h99a, 12'h99b, 12'h99a, 12'h98a, 12'h99b, 12'h99b, 12'h99a, 12'h99a, 12'h88a, 12'h779, 12'h668, 12'h568, 
12'h457, 12'h346, 12'h236, 12'h236, 12'h236, 12'h336, 12'h347, 12'h457, 12'h558, 12'h669, 12'h77a, 12'h99b, 12'haac, 12'hbbd, 12'hcbd, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hbcd, 12'hbbd, 12'hbbd, 12'haad, 12'haac, 12'haac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdef, 12'heee, 12'hede, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hcde, 12'hbbc, 12'h99b, 12'h89a, 12'h89a, 12'h99b, 12'h9ab, 12'h9ab, 12'h89a, 12'h789, 12'h678, 12'h668, 12'h567, 12'h567, 12'h556, 12'h456, 12'h446, 12'h445, 12'h444, 12'h434, 12'h444, 12'h555, 12'h667, 12'h777, 12'h888, 12'h999, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 
12'heed, 12'hedd, 12'hddd, 12'hdcc, 12'hcbb, 12'hbaa, 12'h988, 12'h655, 12'h433, 12'h443, 12'h433, 12'h333, 12'h332, 12'h333, 12'h433, 12'h444, 12'h444, 12'h344, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h333, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h333, 12'h333, 12'h555, 12'h666, 12'h766, 12'h666, 12'h655, 12'h555, 12'h544, 12'h544, 12'h444, 12'h434, 12'h434, 12'h434, 12'h434, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h336, 12'h336, 12'h346, 12'h446, 12'h557, 12'h557, 12'h557, 12'h668, 12'h668, 12'h779, 12'h889, 12'h88a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99a, 12'h99b, 12'h99b, 12'h99a, 12'h88a, 12'h88a, 12'h88a, 12'h879, 12'h779, 12'h668, 12'h668, 12'h668, 12'h568, 
12'h557, 12'h446, 12'h235, 12'h025, 12'h115, 12'h125, 12'h236, 12'h347, 12'h347, 12'h558, 12'h779, 12'h88b, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hbbd, 12'habd, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hedf, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hbbd, 12'h9ab, 12'h89a, 12'h78a, 12'h89a, 12'haab, 12'haab, 12'h89a, 12'h789, 12'h678, 12'h668, 12'h667, 12'h567, 12'h557, 12'h456, 12'h446, 12'h445, 12'h544, 12'h434, 12'h444, 12'h555, 12'h666, 12'h777, 12'h778, 12'h899, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heed, 
12'hedd, 12'hddd, 12'hddd, 12'hdcc, 12'hccb, 12'hbaa, 12'h998, 12'h655, 12'h433, 12'h443, 12'h433, 12'h322, 12'h322, 12'h333, 12'h433, 12'h444, 12'h444, 12'h344, 12'h333, 12'h333, 12'h334, 12'h344, 12'h334, 12'h334, 12'h333, 12'h334, 12'h334, 12'h333, 12'h333, 12'h434, 12'h444, 12'h655, 12'h777, 12'h777, 12'h766, 12'h655, 12'h545, 12'h544, 12'h544, 12'h444, 12'h434, 12'h434, 12'h434, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h336, 12'h336, 12'h446, 12'h446, 12'h446, 12'h557, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h99a, 12'h99b, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'haab, 12'h99b, 12'h99a, 12'h88a, 12'h879, 12'h778, 12'h668, 12'h668, 12'h667, 12'h667, 
12'h567, 12'h457, 12'h336, 12'h235, 12'h225, 12'h335, 12'h346, 12'h447, 12'h347, 12'h447, 12'h669, 12'h88a, 12'h99c, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hbbd, 12'hbbc, 12'haac, 12'haac, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'h99c, 12'haac, 12'haac, 12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heee, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hddf, 12'hdde, 12'hbcd, 12'haac, 12'h89a, 12'h779, 12'h88a, 12'haab, 12'haab, 12'h99a, 12'h789, 12'h678, 12'h668, 12'h667, 12'h567, 12'h557, 12'h456, 12'h456, 12'h445, 12'h545, 12'h445, 12'h445, 12'h555, 12'h666, 12'h777, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'heed, 
12'hedd, 12'hedd, 12'hddd, 12'hdcc, 12'hccb, 12'hbba, 12'h998, 12'h665, 12'h433, 12'h443, 12'h433, 12'h322, 12'h222, 12'h322, 12'h433, 12'h434, 12'h344, 12'h334, 12'h333, 12'h223, 12'h334, 12'h344, 12'h334, 12'h334, 12'h333, 12'h333, 12'h334, 12'h334, 12'h334, 12'h444, 12'h444, 12'h666, 12'h888, 12'h888, 12'h766, 12'h555, 12'h544, 12'h544, 12'h434, 12'h434, 12'h434, 12'h434, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h346, 12'h446, 12'h446, 12'h456, 12'h557, 12'h567, 12'h668, 12'h779, 12'h889, 12'h99a, 12'h99a, 12'haab, 12'haab, 12'haab, 12'hbbb, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbac, 12'haab, 12'h99a, 12'h889, 12'h778, 12'h668, 12'h668, 
12'h667, 12'h557, 12'h456, 12'h446, 12'h446, 12'h557, 12'h668, 12'h668, 12'h457, 12'h337, 12'h558, 12'h77a, 12'h99b, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hbbd, 12'hbbc, 12'haac, 12'haac, 12'h99b, 12'h99b, 12'h99b, 12'h88b, 12'h88a, 12'h78a, 12'h77a, 12'h77a, 12'h88a, 12'h88b, 12'h88b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haac, 12'hbac, 12'hbbc, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hddf, 12'hddf, 12'hdde, 12'hccd, 12'habc, 12'h89b, 12'h669, 12'h78a, 12'haac, 12'habc, 12'h99a, 12'h789, 12'h678, 12'h668, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h555, 12'h555, 12'h545, 12'h545, 12'h556, 12'h666, 12'h777, 12'h778, 12'h889, 12'h9aa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'heee, 12'heed, 12'hedd, 
12'hedd, 12'hedd, 12'hddd, 12'hdcc, 12'hccb, 12'hbaa, 12'h998, 12'h665, 12'h433, 12'h444, 12'h433, 12'h322, 12'h222, 12'h322, 12'h433, 12'h434, 12'h333, 12'h333, 12'h223, 12'h223, 12'h334, 12'h344, 12'h334, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h444, 12'h444, 12'h444, 12'h777, 12'h999, 12'h988, 12'h766, 12'h544, 12'h434, 12'h434, 12'h434, 12'h434, 12'h334, 12'h334, 12'h324, 12'h324, 12'h324, 12'h324, 12'h324, 12'h324, 12'h324, 12'h335, 12'h335, 12'h335, 12'h335, 12'h446, 12'h446, 12'h446, 12'h456, 12'h557, 12'h557, 12'h667, 12'h778, 12'h889, 12'h889, 12'h99a, 12'h99a, 12'haab, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbbc, 12'haab, 12'h99a, 12'h889, 12'h778, 12'h668, 
12'h667, 12'h667, 12'h557, 12'h557, 12'h557, 12'h557, 12'h668, 12'h679, 12'h558, 12'h337, 12'h558, 12'h779, 12'h88b, 12'haac, 12'haac, 12'hbbd, 12'hcce, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hbbc, 12'hbbc, 12'haac, 12'haac, 12'haab, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h78a, 12'h77a, 12'h679, 12'h679, 12'h77a, 12'h77a, 12'h87a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'hbac, 12'hbbc, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 
12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'habc, 12'h89b, 12'h568, 12'h789, 12'haab, 12'habc, 12'h99a, 12'h789, 12'h678, 12'h668, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h555, 12'h655, 12'h555, 12'h555, 12'h556, 12'h666, 12'h777, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heed, 12'hedd, 12'hedd, 
12'hedd, 12'hedd, 12'hddd, 12'hdcc, 12'hcbb, 12'haaa, 12'h988, 12'h665, 12'h543, 12'h544, 12'h443, 12'h322, 12'h221, 12'h322, 12'h434, 12'h434, 12'h333, 12'h333, 12'h223, 12'h223, 12'h333, 12'h344, 12'h334, 12'h333, 12'h333, 12'h333, 12'h334, 12'h334, 12'h444, 12'h444, 12'h444, 12'h777, 12'h999, 12'h999, 12'h766, 12'h544, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h334, 12'h334, 12'h334, 12'h324, 12'h324, 12'h324, 12'h324, 12'h324, 12'h224, 12'h325, 12'h335, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h456, 12'h556, 12'h557, 12'h667, 12'h668, 12'h778, 12'h778, 12'h889, 12'h889, 12'h99a, 12'haab, 12'hbbb, 12'hbbc, 12'hbbc, 12'hcbc, 12'hccd, 12'hccd, 12'hbbc, 12'hbab, 12'h99a, 12'h889, 12'h778, 
12'h667, 12'h557, 12'h446, 12'h446, 12'h457, 12'h557, 12'h778, 12'h779, 12'h558, 12'h226, 12'h447, 12'h669, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hccd, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hede, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hbbc, 12'hbac, 12'haac, 12'haab, 12'haab, 12'haab, 12'ha9b, 12'h99b, 12'h99b, 12'h88b, 12'h88a, 12'h77a, 12'h77a, 12'h779, 12'h77a, 12'h77a, 12'h87a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'haac, 12'hbac, 12'hbbc, 12'hbbd, 12'hcbd, 12'hccd, 12'hccd, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddd, 12'hddd, 12'hdcd, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 
12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hbbd, 12'h99b, 12'h568, 12'h779, 12'haab, 12'haac, 12'h99a, 12'h789, 12'h678, 12'h568, 12'h567, 12'h567, 12'h557, 12'h456, 12'h456, 12'h556, 12'h656, 12'h656, 12'h555, 12'h656, 12'h667, 12'h667, 12'h778, 12'h899, 12'h9aa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddc, 12'hddc, 
12'hddc, 12'hddc, 12'hdcc, 12'hccb, 12'hbba, 12'ha99, 12'h887, 12'h655, 12'h543, 12'h544, 12'h444, 12'h333, 12'h322, 12'h333, 12'h434, 12'h444, 12'h333, 12'h333, 12'h222, 12'h122, 12'h333, 12'h344, 12'h334, 12'h223, 12'h223, 12'h333, 12'h334, 12'h334, 12'h434, 12'h444, 12'h444, 12'h777, 12'h999, 12'h999, 12'h766, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h334, 12'h335, 12'h335, 12'h335, 12'h224, 12'h224, 12'h225, 12'h335, 12'h345, 12'h345, 12'h346, 12'h346, 12'h345, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h445, 12'h556, 12'h556, 12'h778, 12'h889, 12'h99a, 12'h989, 12'h99a, 12'haab, 12'hcbc, 12'hccd, 12'hccd, 12'hcbc, 12'haab, 12'h99a, 12'h889, 
12'h668, 12'h557, 12'h446, 12'h335, 12'h446, 12'h457, 12'h668, 12'h668, 12'h557, 12'h226, 12'h447, 12'h558, 12'h779, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heef, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hcbd, 12'hbbc, 12'hbac, 12'haac, 12'haac, 12'haab, 12'haab, 12'haab, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h99b, 12'ha9b, 12'haac, 12'hbac, 12'hbbd, 12'hcbd, 12'hcbd, 12'hccd, 12'hccd, 12'hdcd, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hddf, 12'hdde, 12'hcde, 12'hbbd, 12'h99b, 12'h568, 12'h779, 12'h9ab, 12'haac, 12'h99a, 12'h789, 12'h678, 12'h668, 12'h567, 12'h567, 12'h456, 12'h456, 12'h556, 12'h556, 12'h656, 12'h656, 12'h555, 12'h656, 12'h667, 12'h667, 12'h778, 12'h899, 12'h99a, 12'haab, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccb, 12'hccb, 12'hccb, 12'hccb, 
12'hccb, 12'hccb, 12'hcbb, 12'hbba, 12'haa9, 12'h988, 12'h776, 12'h654, 12'h443, 12'h544, 12'h544, 12'h433, 12'h322, 12'h333, 12'h444, 12'h444, 12'h334, 12'h333, 12'h223, 12'h122, 12'h333, 12'h344, 12'h334, 12'h223, 12'h223, 12'h333, 12'h333, 12'h333, 12'h334, 12'h434, 12'h433, 12'h777, 12'h999, 12'h999, 12'h766, 12'h534, 12'h434, 12'h434, 12'h544, 12'h545, 12'h545, 12'h545, 12'h445, 12'h445, 12'h445, 12'h435, 12'h435, 12'h335, 12'h335, 12'h235, 12'h224, 12'h224, 12'h235, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h224, 12'h224, 12'h335, 12'h445, 12'h666, 12'h778, 12'h888, 12'h878, 12'h889, 12'ha9a, 12'hbac, 12'hcbc, 12'hccd, 12'hcbc, 12'hbab, 12'haab, 12'h99a, 
12'h778, 12'h667, 12'h446, 12'h335, 12'h335, 12'h346, 12'h557, 12'h668, 12'h447, 12'h226, 12'h337, 12'h548, 12'h669, 12'h77a, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hccd, 12'hccd, 12'hdde, 12'hdde, 12'hdcd, 12'hdcd, 12'hccd, 12'hccd, 12'hccd, 12'hcbd, 12'hbbc, 12'hbbc, 12'hbac, 12'haab, 12'haab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h98b, 12'h99b, 12'h99b, 12'h99b, 12'haac, 12'hbac, 12'hbbd, 12'hcbd, 12'hccd, 12'hccd, 12'hccd, 12'hcbd, 12'hcbd, 12'hcbd, 12'hccd, 12'hdcd, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 
12'hcce, 12'hdde, 12'hdde, 12'hcde, 12'hbbd, 12'h99b, 12'h568, 12'h779, 12'h9ab, 12'haab, 12'h89a, 12'h789, 12'h678, 12'h678, 12'h567, 12'h557, 12'h557, 12'h557, 12'h556, 12'h556, 12'h656, 12'h656, 12'h656, 12'h556, 12'h656, 12'h667, 12'h888, 12'h999, 12'h99a, 12'haab, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'hbaa, 12'haa9, 12'haa9, 12'hbaa, 12'hbaa, 
12'hbaa, 12'hbaa, 12'hbaa, 12'ha99, 12'h887, 12'h766, 12'h655, 12'h543, 12'h433, 12'h544, 12'h544, 12'h433, 12'h333, 12'h333, 12'h444, 12'h444, 12'h444, 12'h334, 12'h223, 12'h223, 12'h333, 12'h344, 12'h334, 12'h223, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h776, 12'h999, 12'h999, 12'h766, 12'h544, 12'h434, 12'h544, 12'h545, 12'h545, 12'h545, 12'h545, 12'h545, 12'h545, 12'h445, 12'h445, 12'h435, 12'h435, 12'h335, 12'h335, 12'h224, 12'h224, 12'h234, 12'h235, 12'h235, 12'h235, 12'h235, 12'h224, 12'h234, 12'h335, 12'h335, 12'h345, 12'h445, 12'h335, 12'h334, 12'h334, 12'h334, 12'h445, 12'h666, 12'h667, 12'h767, 12'h778, 12'h989, 12'ha9b, 12'hbab, 12'hbbc, 12'hbbc, 12'hbbb, 12'haab, 12'haaa, 
12'h989, 12'h778, 12'h556, 12'h335, 12'h225, 12'h225, 12'h446, 12'h557, 12'h447, 12'h336, 12'h337, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99b, 12'haab, 12'haac, 12'haab, 12'h9ab, 12'h9ab, 12'haab, 12'haac, 12'hbbc, 12'hccd, 12'hccd, 12'hccd, 12'hdcd, 12'hdcd, 12'hdce, 12'hdce, 12'hdcd, 12'hccd, 12'hcbd, 12'hbbc, 12'haac, 12'haab, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h98a, 12'h98a, 12'h99b, 12'h99b, 12'haab, 12'hbac, 12'hbbc, 12'hbbd, 12'hcbd, 12'hcbd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hcbc, 12'hcbd, 12'hdcd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbbd, 
12'hbcd, 12'hcde, 12'hdde, 12'hcde, 12'hbbd, 12'h9ab, 12'h779, 12'h789, 12'h99b, 12'h9ab, 12'h89a, 12'h789, 12'h678, 12'h668, 12'h567, 12'h567, 12'h457, 12'h457, 12'h557, 12'h556, 12'h656, 12'h656, 12'h656, 12'h556, 12'h656, 12'h667, 12'h778, 12'h889, 12'h99a, 12'haab, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hedd, 12'hdcc, 12'hbbb, 12'haa9, 12'h988, 12'h887, 12'h887, 12'h987, 12'h988, 
12'h998, 12'h998, 12'h988, 12'h887, 12'h765, 12'h543, 12'h432, 12'h421, 12'h422, 12'h443, 12'h444, 12'h433, 12'h333, 12'h333, 12'h444, 12'h444, 12'h444, 12'h344, 12'h223, 12'h223, 12'h333, 12'h444, 12'h334, 12'h223, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h222, 12'h666, 12'h999, 12'h999, 12'h767, 12'h545, 12'h545, 12'h656, 12'h656, 12'h666, 12'h667, 12'h667, 12'h667, 12'h667, 12'h657, 12'h556, 12'h446, 12'h446, 12'h335, 12'h335, 12'h225, 12'h225, 12'h235, 12'h235, 12'h235, 12'h235, 12'h335, 12'h335, 12'h335, 12'h445, 12'h446, 12'h446, 12'h446, 12'h445, 12'h335, 12'h335, 12'h335, 12'h446, 12'h556, 12'h667, 12'h668, 12'h878, 12'h99a, 12'hbac, 12'hbbc, 12'hcbc, 12'hbbc, 12'hbab, 12'haab, 12'ha9a, 
12'h989, 12'h778, 12'h557, 12'h446, 12'h335, 12'h335, 12'h447, 12'h557, 12'h447, 12'h226, 12'h337, 12'h447, 12'h558, 12'h769, 12'h77a, 12'h88a, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'habc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hccd, 12'hccd, 12'hdce, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'hbbc, 12'haac, 12'haab, 12'haab, 12'h99b, 12'h99a, 12'h98a, 12'h99a, 12'h99a, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h769, 12'h779, 12'h779, 12'h88a, 12'h99a, 12'h99b, 12'h99b, 12'h99b, 12'ha9b, 12'haab, 12'haac, 12'hbac, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdcd, 12'hccc, 
12'hcbc, 12'hccd, 12'hddd, 12'hddd, 12'hccd, 12'haab, 12'h88a, 12'h889, 12'h89a, 12'h89a, 12'h88a, 12'h889, 12'h779, 12'h668, 12'h568, 12'h568, 12'h467, 12'h457, 12'h457, 12'h557, 12'h656, 12'h556, 12'h556, 12'h556, 12'h656, 12'h667, 12'h777, 12'h888, 12'h99a, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbba, 12'ha99, 12'h887, 12'h765, 12'h765, 12'h766, 12'h766, 
12'h777, 12'h877, 12'h776, 12'h766, 12'h655, 12'h443, 12'h433, 12'h322, 12'h433, 12'h433, 12'h444, 12'h433, 12'h433, 12'h433, 12'h444, 12'h444, 12'h444, 12'h444, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h334, 12'h333, 12'h333, 12'h334, 12'h334, 12'h323, 12'h313, 12'h767, 12'h999, 12'ha9a, 12'h778, 12'h656, 12'h656, 12'h767, 12'h778, 12'h889, 12'h889, 12'h98a, 12'h88a, 12'h88a, 12'h779, 12'h668, 12'h558, 12'h447, 12'h346, 12'h236, 12'h236, 12'h236, 12'h236, 12'h236, 12'h346, 12'h446, 12'h446, 12'h557, 12'h557, 12'h557, 12'h557, 12'h557, 12'h447, 12'h446, 12'h446, 12'h447, 12'h447, 12'h457, 12'h558, 12'h668, 12'h769, 12'h98a, 12'hbac, 12'hdcd, 12'hdce, 12'hdcd, 12'hccd, 12'haab, 12'h99a, 12'h98a, 
12'h889, 12'h778, 12'h667, 12'h546, 12'h446, 12'h446, 12'h557, 12'h557, 12'h447, 12'h226, 12'h337, 12'h548, 12'h669, 12'h77a, 12'h88a, 12'h88b, 12'h99b, 12'h99c, 12'haac, 12'hbad, 12'hbbd, 12'hbbd, 12'hbbd, 12'habc, 12'haac, 12'haac, 12'haac, 12'haac, 12'hbbc, 12'hccd, 12'hdce, 12'hddf, 12'hedf, 12'hdde, 12'hccd, 12'hbbd, 12'hbac, 12'haab, 12'haab, 12'ha9b, 12'h99a, 12'h88a, 12'h88a, 12'h88a, 12'h779, 12'h768, 12'h658, 12'h547, 12'h447, 12'h557, 12'h658, 12'h668, 12'h779, 12'h779, 12'h779, 12'h779, 12'h88a, 12'h98a, 12'h99b, 12'haac, 12'hbbc, 12'hbbc, 12'hbbc, 12'haac, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'hede, 12'hede, 12'heee, 12'heee, 12'hdde, 12'hccd, 
12'hcbc, 12'hccd, 12'hccd, 12'hccd, 12'hccc, 12'hbbb, 12'h99a, 12'h889, 12'h889, 12'h889, 12'h889, 12'h889, 12'h779, 12'h668, 12'h668, 12'h568, 12'h568, 12'h357, 12'h457, 12'h557, 12'h657, 12'h556, 12'h556, 12'h656, 12'h656, 12'h667, 12'h777, 12'h888, 12'h99a, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccc, 12'hbba, 12'h999, 12'h877, 12'h665, 12'h654, 12'h545, 12'h545, 
12'h545, 12'h545, 12'h545, 12'h545, 12'h544, 12'h434, 12'h434, 12'h433, 12'h333, 12'h433, 12'h434, 12'h433, 12'h433, 12'h434, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h434, 12'h323, 12'h434, 12'h434, 12'h434, 12'h324, 12'h323, 12'h424, 12'h434, 12'h424, 12'h313, 12'h767, 12'ha9a, 12'haaa, 12'h878, 12'h767, 12'h768, 12'h879, 12'h88a, 12'h99b, 12'haab, 12'haac, 12'haac, 12'h9ab, 12'h89b, 12'h78a, 12'h669, 12'h458, 12'h247, 12'h136, 12'h136, 12'h236, 12'h236, 12'h336, 12'h447, 12'h557, 12'h557, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h558, 12'h558, 12'h558, 12'h558, 12'h558, 12'h558, 12'h669, 12'h669, 12'h879, 12'h98b, 12'hcbc, 12'hede, 12'hede, 12'hdde, 12'hccd, 12'hbab, 12'h99a, 12'h99a, 
12'h98a, 12'h889, 12'h668, 12'h657, 12'h657, 12'h557, 12'h668, 12'h668, 12'h547, 12'h336, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99b, 12'h99c, 12'haac, 12'hbbd, 12'hbbd, 12'hcbd, 12'hcbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'hcbd, 12'hcce, 12'hdde, 12'hddf, 12'hdde, 12'hcce, 12'hcbd, 12'hbbc, 12'haac, 12'ha9b, 12'h99a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h779, 12'h668, 12'h557, 12'h436, 12'h326, 12'h436, 12'h447, 12'h547, 12'h557, 12'h557, 12'h447, 12'h557, 12'h668, 12'h779, 12'h98a, 12'ha9b, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'habd, 12'hbbd, 12'hccd, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hede, 12'hddd, 
12'hccd, 12'hcbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'haab, 12'h889, 12'h778, 12'h779, 12'h779, 12'h889, 12'h789, 12'h779, 12'h668, 12'h568, 12'h568, 12'h458, 12'h357, 12'h457, 12'h557, 12'h667, 12'h657, 12'h657, 12'h656, 12'h666, 12'h667, 12'h777, 12'h888, 12'ha9a, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccc, 12'hbba, 12'h998, 12'h876, 12'h655, 12'h544, 12'h434, 12'h334, 
12'h324, 12'h334, 12'h334, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h334, 12'h334, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h444, 12'h544, 12'h544, 12'h434, 12'h323, 12'h423, 12'h444, 12'h434, 12'h424, 12'h323, 12'h424, 12'h435, 12'h435, 12'h324, 12'h767, 12'ha9a, 12'haab, 12'h989, 12'h879, 12'h879, 12'h98a, 12'h99b, 12'haab, 12'hbac, 12'hbbc, 12'hbbc, 12'haac, 12'h99b, 12'h78a, 12'h679, 12'h458, 12'h247, 12'h137, 12'h137, 12'h237, 12'h337, 12'h447, 12'h557, 12'h668, 12'h668, 12'h779, 12'h779, 12'h889, 12'h889, 12'h889, 12'h88a, 12'h88a, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h99b, 12'hbac, 12'hcbd, 12'hdde, 12'hede, 12'hede, 12'hdde, 12'hcbd, 12'hbbc, 12'haab, 
12'haab, 12'h99a, 12'h879, 12'h778, 12'h778, 12'h768, 12'h668, 12'h668, 12'h558, 12'h558, 12'h558, 12'h558, 12'h669, 12'h87a, 12'h99b, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hbbc, 12'haac, 12'h99b, 12'h88a, 12'h88a, 12'h88a, 12'h98a, 12'h99a, 12'h88a, 12'h779, 12'h668, 12'h547, 12'h436, 12'h447, 12'h447, 12'h447, 12'h447, 12'h437, 12'h336, 12'h447, 12'h658, 12'h779, 12'h88a, 12'h99b, 12'ha9b, 12'ha9b, 12'haab, 12'haac, 12'habc, 12'haac, 12'haac, 12'hbbd, 12'hbcd, 12'hccd, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'hdde, 
12'hdcd, 12'hbbb, 12'haaa, 12'haaa, 12'haab, 12'h99a, 12'h878, 12'h778, 12'h778, 12'h778, 12'h779, 12'h779, 12'h678, 12'h568, 12'h568, 12'h568, 12'h568, 12'h457, 12'h457, 12'h557, 12'h667, 12'h657, 12'h657, 12'h656, 12'h667, 12'h667, 12'h777, 12'h889, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccc, 12'hbaa, 12'h998, 12'h876, 12'h654, 12'h433, 12'h333, 12'h324, 
12'h324, 12'h334, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h334, 12'h333, 12'h333, 12'h333, 12'h323, 12'h323, 12'h323, 12'h433, 12'h434, 12'h444, 12'h434, 12'h433, 12'h323, 12'h323, 12'h434, 12'h434, 12'h424, 12'h324, 12'h434, 12'h435, 12'h435, 12'h434, 12'h767, 12'ha9a, 12'haab, 12'h99a, 12'h98a, 12'h98a, 12'h99a, 12'ha9b, 12'haab, 12'haac, 12'hbbc, 12'haac, 12'haac, 12'h99b, 12'h88a, 12'h679, 12'h568, 12'h358, 12'h347, 12'h347, 12'h347, 12'h457, 12'h558, 12'h568, 12'h668, 12'h779, 12'h889, 12'h88a, 12'h99a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'haac, 12'hbac, 12'hcbd, 12'hccd, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'hcbc, 
12'hbbc, 12'haab, 12'h99a, 12'h889, 12'h889, 12'h779, 12'h668, 12'h668, 12'h668, 12'h669, 12'h669, 12'h558, 12'h669, 12'h88a, 12'h99b, 12'hbbd, 12'hcce, 12'hcce, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hbbd, 12'haac, 12'haac, 12'hbbd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hdce, 12'hccd, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h98a, 12'h99a, 12'h99b, 12'h99b, 12'h99a, 12'h879, 12'h779, 12'h658, 12'h547, 12'h547, 12'h547, 12'h447, 12'h447, 12'h437, 12'h336, 12'h447, 12'h668, 12'h779, 12'h88a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'hede, 
12'hccd, 12'haab, 12'h989, 12'h989, 12'h99a, 12'h889, 12'h778, 12'h667, 12'h668, 12'h668, 12'h778, 12'h778, 12'h678, 12'h568, 12'h568, 12'h568, 12'h568, 12'h457, 12'h457, 12'h557, 12'h667, 12'h657, 12'h657, 12'h657, 12'h667, 12'h767, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hccc, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccc, 12'hbaa, 12'h998, 12'h776, 12'h654, 12'h433, 12'h333, 12'h324, 
12'h334, 12'h334, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h444, 12'h434, 12'h434, 12'h434, 12'h433, 12'h433, 12'h433, 12'h333, 12'h333, 12'h433, 12'h433, 12'h433, 12'h433, 12'h433, 12'h323, 12'h433, 12'h434, 12'h434, 12'h324, 12'h323, 12'h424, 12'h435, 12'h435, 12'h435, 12'h767, 12'h999, 12'ha9a, 12'ha9a, 12'h99a, 12'h99a, 12'h99a, 12'h99b, 12'h99b, 12'haab, 12'haab, 12'haac, 12'h9ac, 12'h99b, 12'h88a, 12'h77a, 12'h679, 12'h569, 12'h568, 12'h568, 12'h568, 12'h568, 12'h668, 12'h669, 12'h779, 12'h779, 12'h88a, 12'h98a, 12'h99b, 12'ha9b, 12'haab, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'habd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hcbd, 12'hccd, 12'hccd, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdcd, 
12'hcbc, 12'hbbc, 12'haab, 12'h99a, 12'h99a, 12'h889, 12'h678, 12'h568, 12'h668, 12'h779, 12'h779, 12'h669, 12'h779, 12'h99b, 12'haac, 12'hcbd, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hcce, 12'hccd, 12'hcce, 12'hcce, 12'hbbd, 12'hbbc, 12'hbbc, 12'hccd, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hbbc, 12'ha9b, 12'h99b, 12'h99b, 12'haab, 12'haab, 12'haab, 12'h99b, 12'h88a, 12'h889, 12'h779, 12'h668, 12'h668, 12'h668, 12'h558, 12'h547, 12'h447, 12'h447, 12'h557, 12'h668, 12'h879, 12'h88a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'h9ac, 12'h99b, 12'h99b, 12'haac, 12'hbbc, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'hdde, 
12'hccd, 12'h99a, 12'h878, 12'h888, 12'h889, 12'h878, 12'h667, 12'h667, 12'h667, 12'h667, 12'h668, 12'h678, 12'h668, 12'h568, 12'h668, 12'h668, 12'h568, 12'h568, 12'h557, 12'h557, 12'h667, 12'h657, 12'h557, 12'h657, 12'h667, 12'h767, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hccd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hcbb, 12'haaa, 12'h998, 12'h776, 12'h654, 12'h544, 12'h434, 12'h434, 
12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h444, 12'h444, 12'h444, 12'h444, 12'h544, 12'h544, 12'h544, 12'h444, 12'h444, 12'h434, 12'h434, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h434, 12'h434, 12'h323, 12'h323, 12'h424, 12'h434, 12'h434, 12'h434, 12'h656, 12'h889, 12'h99a, 12'ha9a, 12'ha9b, 12'h99a, 12'h98a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h89b, 12'h89b, 12'h88b, 12'h88a, 12'h78a, 12'h78a, 12'h77a, 12'h77a, 12'h77a, 12'h779, 12'h679, 12'h779, 12'h779, 12'h879, 12'h88a, 12'h88a, 12'h99a, 12'h99b, 12'haab, 12'haac, 12'haac, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hcbd, 12'hcbd, 12'hcbd, 12'hcbd, 12'hcbd, 12'hccd, 12'hdde, 12'hdde, 12'hdde, 
12'hccd, 12'hbbc, 12'haab, 12'haab, 12'h99a, 12'h88a, 12'h678, 12'h668, 12'h668, 12'h779, 12'h779, 12'h779, 12'h77a, 12'h99c, 12'hbbd, 12'hcce, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hbbd, 12'hbbc, 12'hbbd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hbbd, 12'hbac, 12'haac, 12'haac, 12'haac, 12'hbac, 12'hbac, 12'haac, 12'ha9b, 12'h99b, 12'h98a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h779, 12'h879, 12'h98a, 12'h99b, 12'haab, 12'haac, 12'haac, 12'haab, 12'haab, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'haac, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'hddd, 12'hdcd, 12'hccd, 
12'hbbc, 12'h989, 12'h778, 12'h778, 12'h889, 12'h778, 12'h667, 12'h667, 12'h557, 12'h567, 12'h667, 12'h668, 12'h668, 12'h567, 12'h568, 12'h668, 12'h568, 12'h568, 12'h568, 12'h557, 12'h557, 12'h557, 12'h657, 12'h667, 12'h667, 12'h778, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hedd, 12'hdcc, 12'hbbb, 12'haa9, 12'h988, 12'h876, 12'h665, 12'h655, 12'h555, 12'h545, 
12'h545, 12'h545, 12'h444, 12'h434, 12'h434, 12'h434, 12'h444, 12'h544, 12'h545, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h555, 12'h444, 12'h444, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h323, 12'h323, 12'h323, 12'h424, 12'h434, 12'h434, 12'h656, 12'h778, 12'h989, 12'ha9b, 12'haab, 12'ha9b, 12'h98a, 12'h88a, 12'h779, 12'h779, 12'h78a, 12'h88a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 12'h88b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h98a, 12'h99b, 12'h99b, 12'ha9b, 12'haac, 12'haac, 12'hbac, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hbbd, 12'hbac, 12'hbac, 12'hbac, 12'hbac, 12'hbbc, 12'hcbd, 12'hbbc, 
12'hbbc, 12'haab, 12'haab, 12'h99a, 12'h88a, 12'h889, 12'h779, 12'h668, 12'h669, 12'h779, 12'h779, 12'h77a, 12'h88b, 12'haac, 12'hbbd, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hcce, 12'hccd, 12'hbbd, 12'haac, 12'haac, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hcbd, 12'hbbd, 12'hbbc, 12'hbac, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'hbbc, 12'hbbd, 12'hcbd, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'hccd, 12'hbbc, 12'hbbb, 12'haab, 
12'h99a, 12'h878, 12'h767, 12'h778, 12'h889, 12'h778, 12'h667, 12'h667, 12'h556, 12'h556, 12'h557, 12'h567, 12'h567, 12'h567, 12'h568, 12'h668, 12'h668, 12'h568, 12'h568, 12'h557, 12'h557, 12'h557, 12'h657, 12'h667, 12'h667, 12'h768, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haa9, 12'h998, 12'h887, 12'h776, 12'h766, 12'h766, 12'h666, 
12'h656, 12'h656, 12'h555, 12'h545, 12'h545, 12'h545, 12'h555, 12'h555, 12'h555, 12'h655, 12'h655, 12'h655, 12'h655, 12'h555, 12'h555, 12'h555, 12'h544, 12'h444, 12'h444, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h423, 12'h324, 12'h323, 12'h323, 12'h424, 12'h434, 12'h545, 12'h667, 12'h878, 12'ha9a, 12'haab, 12'haab, 12'h99a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'h99c, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h98b, 12'h99b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbc, 12'hbac, 12'hbac, 12'ha9b, 12'h98a, 12'h88a, 12'h99a, 12'h99b, 12'h99b, 
12'h99a, 12'h99a, 12'h99a, 12'h88a, 12'h789, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h779, 12'h88a, 12'h99b, 12'hbbd, 12'hcce, 12'hdce, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hcce, 12'hcbd, 12'haac, 12'h99b, 12'h99b, 12'haac, 12'hcbd, 12'hdde, 12'hedf, 12'hddf, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hedf, 12'hdde, 12'hccd, 12'hbbc, 12'h99a, 12'h99a, 12'h98a, 
12'h889, 12'h778, 12'h667, 12'h778, 12'h888, 12'h778, 12'h767, 12'h667, 12'h556, 12'h446, 12'h456, 12'h557, 12'h557, 12'h567, 12'h567, 12'h668, 12'h678, 12'h678, 12'h668, 12'h567, 12'h557, 12'h557, 12'h657, 12'h667, 12'h668, 12'h668, 12'h778, 12'h889, 12'haaa, 12'hbbb, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbba, 12'haa9, 12'h999, 12'h988, 12'h887, 12'h887, 12'h878, 12'h777, 
12'h777, 12'h767, 12'h666, 12'h666, 12'h656, 12'h656, 12'h656, 12'h656, 12'h666, 12'h666, 12'h666, 12'h666, 12'h655, 12'h655, 12'h655, 12'h555, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h434, 12'h434, 12'h433, 12'h423, 12'h323, 12'h323, 12'h324, 12'h434, 12'h434, 12'h546, 12'h767, 12'h99a, 12'haab, 12'haab, 12'h99a, 12'h99a, 12'h88a, 12'h88a, 12'h99b, 12'h99c, 12'haac, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h88a, 12'h88a, 12'h98b, 12'h99b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haac, 12'haad, 12'haad, 12'hbad, 12'hbac, 12'hbac, 12'haac, 12'h99b, 12'h87a, 12'h668, 12'h769, 12'h779, 12'h779, 
12'h889, 12'h889, 12'h88a, 12'h779, 12'h679, 12'h668, 12'h779, 12'h88a, 12'h88a, 12'h779, 12'h77a, 12'h88a, 12'h99b, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hcce, 12'hbbd, 12'haac, 12'h88a, 12'h88a, 12'h99b, 12'hbac, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'hbbd, 12'haac, 12'hbac, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hccd, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hbbc, 12'h99a, 12'h779, 12'h778, 12'h889, 
12'h889, 12'h767, 12'h667, 12'h778, 12'h878, 12'h778, 12'h767, 12'h667, 12'h556, 12'h446, 12'h446, 12'h456, 12'h457, 12'h557, 12'h567, 12'h567, 12'h668, 12'h678, 12'h668, 12'h568, 12'h557, 12'h557, 12'h668, 12'h668, 12'h678, 12'h778, 12'h778, 12'h999, 12'haab, 12'hbbc, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'hbaa, 12'haa9, 12'ha99, 12'h999, 12'h999, 12'h999, 12'h989, 
12'h888, 12'h888, 12'h888, 12'h877, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h766, 12'h666, 12'h665, 12'h655, 12'h555, 12'h544, 12'h444, 12'h433, 12'h433, 12'h443, 12'h444, 12'h433, 12'h433, 12'h434, 12'h433, 12'h434, 12'h434, 12'h424, 12'h434, 12'h434, 12'h434, 12'h545, 12'h656, 12'h778, 12'h88a, 12'h88a, 12'h889, 12'h88a, 12'h88a, 12'h88a, 12'h99b, 12'h9ac, 12'haac, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'ha9b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'ha9c, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 12'hbad, 12'hbad, 12'hbac, 12'haac, 12'h99b, 12'h779, 12'h668, 12'h668, 12'h668, 12'h769, 
12'h779, 12'h779, 12'h779, 12'h668, 12'h568, 12'h568, 12'h779, 12'h89a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h99c, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hcce, 12'hbbd, 12'haab, 12'h87a, 12'h779, 12'h99b, 12'haac, 12'hccd, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'hbbd, 12'haac, 12'haac, 12'hbac, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'haab, 12'h889, 12'h657, 12'h657, 12'h778, 
12'h889, 12'h667, 12'h657, 12'h767, 12'h778, 12'h778, 12'h667, 12'h557, 12'h456, 12'h446, 12'h446, 12'h456, 12'h457, 12'h557, 12'h567, 12'h567, 12'h567, 12'h568, 12'h668, 12'h668, 12'h568, 12'h668, 12'h668, 12'h668, 12'h778, 12'h778, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hcbb, 12'hbbb, 12'hbaa, 12'haa9, 12'haa9, 12'haa9, 12'ha99, 
12'h999, 12'h999, 12'h999, 12'h999, 12'h988, 12'h988, 12'h988, 12'h888, 12'h888, 12'h888, 12'h887, 12'h877, 12'h777, 12'h766, 12'h666, 12'h655, 12'h554, 12'h544, 12'h544, 12'h444, 12'h443, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h545, 12'h557, 12'h658, 12'h668, 12'h668, 12'h779, 12'h77a, 12'h88a, 12'h99b, 12'h99c, 12'haac, 12'haad, 12'habd, 12'habd, 12'habd, 12'hbbd, 12'hbbe, 12'hbce, 12'hbce, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 12'haad, 12'hbad, 12'hbad, 12'hbac, 12'haac, 12'h99b, 12'h779, 12'h658, 12'h668, 12'h668, 12'h668, 
12'h669, 12'h669, 12'h668, 12'h558, 12'h558, 12'h558, 12'h78a, 12'h99b, 12'h89b, 12'h88a, 12'h88b, 12'h88b, 12'h99c, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hdde, 12'hcce, 12'hccd, 12'haac, 12'h88a, 12'h87a, 12'h99b, 12'hbac, 12'hccd, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdce, 12'hccd, 12'hbbd, 12'hbbc, 12'hbac, 12'hbac, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdce, 12'hcce, 12'hccd, 12'hcbd, 12'haac, 12'h98a, 12'h768, 12'h446, 12'h557, 12'h879, 
12'h889, 12'h667, 12'h556, 12'h667, 12'h778, 12'h767, 12'h667, 12'h557, 12'h456, 12'h446, 12'h446, 12'h456, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h568, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h778, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hccb, 12'hbbb, 12'hbaa, 12'haaa, 12'haaa, 12'haaa, 
12'ha99, 12'ha99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h998, 12'h888, 12'h888, 12'h887, 12'h777, 12'h776, 12'h666, 12'h665, 12'h665, 12'h655, 12'h555, 12'h544, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h444, 12'h444, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h436, 12'h447, 12'h547, 12'h558, 12'h668, 12'h779, 12'h78a, 12'h88a, 12'h89b, 12'h99c, 12'h99c, 12'h9ac, 12'h9ac, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbac, 12'ha9c, 12'h98b, 12'h77a, 12'h669, 12'h769, 12'h779, 12'h779, 
12'h669, 12'h668, 12'h558, 12'h457, 12'h447, 12'h558, 12'h78a, 12'h99b, 12'h99b, 12'h88b, 12'h88b, 12'h89b, 12'h99c, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdce, 12'hccd, 12'hbbc, 12'h99b, 12'h99b, 12'hbbc, 12'hccd, 12'hdce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hcce, 12'hccd, 12'hcbd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdce, 12'hcce, 12'hbbd, 12'hbbc, 12'haab, 12'h99a, 12'h779, 12'h658, 12'h446, 12'h657, 12'h889, 
12'h889, 12'h667, 12'h546, 12'h556, 12'h667, 12'h667, 12'h667, 12'h557, 12'h456, 12'h446, 12'h456, 12'h557, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h778, 12'h779, 12'h789, 12'h889, 12'h99a, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hdcc, 12'hccb, 12'hbbb, 12'hbaa, 12'haaa, 12'haaa, 
12'ha99, 12'h999, 12'h999, 12'h999, 12'h999, 12'h998, 12'h998, 12'h998, 12'h998, 12'h998, 12'h998, 12'h888, 12'h888, 12'h887, 12'h877, 12'h777, 12'h777, 12'h777, 12'h776, 12'h666, 12'h555, 12'h433, 12'h433, 12'h433, 12'h433, 12'h444, 12'h444, 12'h444, 12'h444, 12'h434, 12'h434, 12'h434, 12'h434, 12'h434, 12'h435, 12'h436, 12'h447, 12'h547, 12'h558, 12'h669, 12'h679, 12'h77a, 12'h78a, 12'h78b, 12'h88b, 12'h89b, 12'h89c, 12'h89c, 12'h99c, 12'h9ac, 12'haad, 12'habd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcbd, 12'hcbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h87a, 12'h77a, 12'h87a, 12'h88a, 12'h779, 
12'h669, 12'h558, 12'h447, 12'h347, 12'h447, 12'h558, 12'h77a, 12'h89b, 12'h89b, 12'h88b, 12'h88b, 12'h99b, 12'haac, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdce, 12'hbbd, 12'haac, 12'haac, 12'hccd, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hcce, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h768, 12'h668, 12'h557, 12'h668, 12'h879, 
12'h879, 12'h657, 12'h446, 12'h556, 12'h667, 12'h667, 12'h667, 12'h557, 12'h456, 12'h446, 12'h456, 12'h557, 12'h567, 12'h567, 12'h567, 12'h567, 12'h567, 12'h568, 12'h678, 12'h668, 12'h668, 12'h668, 12'h668, 12'h778, 12'h779, 12'h789, 12'h89a, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hdcc, 12'hccb, 12'hbbb, 12'hbba, 12'haaa, 
12'haaa, 12'haaa, 12'haaa, 12'haa9, 12'haa9, 12'haa9, 12'haa9, 12'haa9, 12'haa9, 12'haaa, 12'haaa, 12'haa9, 12'haa9, 12'h999, 12'h999, 12'h999, 12'h998, 12'h998, 12'h998, 12'h887, 12'h766, 12'h544, 12'h443, 12'h433, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h434, 12'h433, 12'h433, 12'h434, 12'h434, 12'h335, 12'h336, 12'h437, 12'h447, 12'h558, 12'h568, 12'h669, 12'h77a, 12'h78a, 12'h88b, 12'h89b, 12'h89c, 12'h89c, 12'h99c, 12'h9ad, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbad, 12'hbad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'h99b, 12'h88b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h779, 
12'h669, 12'h458, 12'h337, 12'h237, 12'h447, 12'h558, 12'h77a, 12'h89b, 12'h88b, 12'h78a, 12'h88b, 12'h99c, 12'haac, 12'hbbd, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hccd, 12'hbbd, 12'hbbd, 12'hdce, 12'hdde, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hccd, 12'hcbd, 12'hcbd, 12'hcbd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hcce, 12'hbbc, 12'h99b, 12'h879, 12'h768, 12'h668, 12'h668, 12'h668, 12'h768, 12'h778, 
12'h778, 12'h557, 12'h446, 12'h446, 12'h557, 12'h557, 12'h557, 12'h557, 12'h456, 12'h446, 12'h557, 12'h567, 12'h567, 12'h667, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h679, 12'h669, 12'h668, 12'h679, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hddc, 12'hccc, 12'hccc, 12'hccc, 
12'hcbb, 12'hcbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hcbb, 12'hcbb, 12'hcbb, 12'hcbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbba, 12'hbba, 12'hbba, 12'haaa, 12'haa9, 12'h887, 12'h655, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h433, 12'h323, 12'h323, 12'h433, 12'h434, 12'h325, 12'h226, 12'h336, 12'h337, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h89c, 12'h9ac, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'haad, 12'hbad, 12'hbad, 12'hbad, 12'haad, 12'haad, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haad, 12'haad, 12'hbbd, 12'hbbd, 12'haac, 12'h98b, 12'h88a, 12'h88a, 12'h88b, 12'h88a, 12'h88a, 12'h779, 
12'h558, 12'h447, 12'h116, 12'h126, 12'h448, 12'h569, 12'h77a, 12'h88b, 12'h88b, 12'h77a, 12'h88b, 12'h99c, 12'habd, 12'hcce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hdce, 12'hdce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hbbd, 12'h99b, 12'h879, 12'h769, 12'h768, 12'h779, 12'h879, 12'h879, 12'h779, 
12'h768, 12'h557, 12'h446, 12'h446, 12'h556, 12'h556, 12'h556, 12'h556, 12'h446, 12'h446, 12'h557, 12'h567, 12'h667, 12'h667, 12'h567, 12'h567, 12'h567, 12'h678, 12'h678, 12'h678, 12'h679, 12'h669, 12'h668, 12'h678, 12'h779, 12'h88a, 12'h99a, 12'haab, 12'hccc, 12'hcdd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'hedd, 12'hddd, 12'hddd, 12'hddd, 
12'hddd, 12'hddc, 12'hddc, 12'hdcc, 12'hdcc, 12'hdcc, 12'hddc, 12'hddc, 12'hddc, 12'hddc, 12'hddc, 12'hddc, 12'hddc, 12'hdcc, 12'hccc, 12'hccc, 12'hccc, 12'hccb, 12'hccb, 12'hbba, 12'h999, 12'h766, 12'h554, 12'h544, 12'h544, 12'h434, 12'h444, 12'h444, 12'h444, 12'h333, 12'h212, 12'h322, 12'h434, 12'h434, 12'h325, 12'h216, 12'h226, 12'h226, 12'h347, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99c, 12'h9ad, 12'haad, 12'habd, 12'habe, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbad, 12'hbad, 12'hbad, 12'hbad, 12'hbad, 12'hbad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'h99b, 12'h99b, 12'ha9c, 12'haac, 12'haac, 12'h99b, 12'h88b, 
12'h77a, 12'h669, 12'h458, 12'h448, 12'h458, 12'h569, 12'h67a, 12'h78a, 12'h78a, 12'h77a, 12'h88b, 12'h99c, 12'hbbd, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hddf, 12'hedf, 12'hdce, 12'haac, 12'h99b, 12'h88a, 12'h889, 12'h88a, 12'h98a, 12'h98a, 12'h889, 
12'h778, 12'h667, 12'h556, 12'h556, 12'h557, 12'h557, 12'h557, 12'h556, 12'h446, 12'h446, 12'h556, 12'h567, 12'h567, 12'h567, 12'h567, 12'h557, 12'h567, 12'h668, 12'h678, 12'h678, 12'h679, 12'h669, 12'h668, 12'h679, 12'h779, 12'h88a, 12'h99a, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'heee, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heee, 12'heed, 12'heed, 12'heed, 12'heed, 12'hedd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddc, 12'hdcc, 12'hddc, 12'hddc, 12'hdcc, 12'hccb, 12'haa9, 12'h776, 12'h655, 12'h554, 12'h544, 12'h444, 12'h444, 12'h444, 12'h444, 12'h433, 12'h222, 12'h323, 12'h444, 12'h445, 12'h435, 12'h226, 12'h226, 12'h337, 12'h347, 12'h448, 12'h559, 12'h669, 12'h77a, 12'h78b, 12'h89c, 12'h99c, 12'h9ad, 12'haad, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbce, 12'hbbe, 12'hbbd, 12'hbac, 12'haac, 12'haac, 12'hbbd, 12'hccd, 12'hbbd, 12'hbbd, 12'haac, 
12'h99b, 12'h89b, 12'h77a, 12'h669, 12'h569, 12'h569, 12'h669, 12'h67a, 12'h77a, 12'h78b, 12'h89b, 12'h9ac, 12'hbbd, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hbbd, 12'hcbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'hdde, 12'hbbd, 12'ha9b, 12'h98a, 12'h88a, 12'h98a, 12'h99a, 12'h99a, 12'h889, 
12'h778, 12'h768, 12'h668, 12'h668, 12'h778, 12'h778, 12'h778, 12'h667, 12'h556, 12'h446, 12'h456, 12'h557, 12'h567, 12'h667, 12'h567, 12'h557, 12'h567, 12'h668, 12'h678, 12'h678, 12'h669, 12'h669, 12'h669, 12'h779, 12'h789, 12'h88a, 12'h99b, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hffe, 12'hffe, 12'hffe, 12'hfee, 12'hfee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heed, 12'hedd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hbaa, 12'h887, 12'h666, 12'h555, 12'h544, 12'h444, 12'h443, 12'h444, 12'h444, 12'h433, 12'h322, 12'h333, 12'h544, 12'h545, 12'h446, 12'h336, 12'h337, 12'h337, 12'h347, 12'h348, 12'h458, 12'h569, 12'h66a, 12'h77b, 12'h78b, 12'h89c, 12'h99c, 12'h9ad, 12'haae, 12'habe, 12'hbbe, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbbe, 12'hbbd, 12'hbad, 12'hbbd, 12'hbbd, 12'hcce, 12'hdce, 12'hcce, 12'hbcd, 12'hbbd, 
12'haac, 12'h99b, 12'h78a, 12'h679, 12'h669, 12'h569, 12'h569, 12'h67a, 12'h77a, 12'h88b, 12'h99c, 12'haad, 12'hbbd, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hdde, 12'hcbd, 12'hbac, 12'h99b, 12'h98a, 12'h88a, 12'h88a, 12'h879, 12'h779, 
12'h779, 12'h889, 12'h88a, 12'h99a, 12'ha9b, 12'haab, 12'haab, 12'h99a, 12'h668, 12'h446, 12'h346, 12'h456, 12'h567, 12'h668, 12'h667, 12'h557, 12'h567, 12'h667, 12'h678, 12'h668, 12'h668, 12'h669, 12'h679, 12'h779, 12'h889, 12'h88a, 12'h9ab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'heee, 12'heee, 12'heed, 12'heed, 12'heed, 12'heed, 12'heed, 12'heed, 12'hddc, 12'hbbb, 12'h988, 12'h776, 12'h655, 12'h544, 12'h544, 12'h443, 12'h433, 12'h433, 12'h433, 12'h433, 12'h434, 12'h544, 12'h545, 12'h336, 12'h336, 12'h226, 12'h237, 12'h337, 12'h348, 12'h448, 12'h559, 12'h56a, 12'h67a, 12'h78b, 12'h78c, 12'h89c, 12'h99d, 12'h9ad, 12'haad, 12'haad, 12'haae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 
12'haac, 12'h99b, 12'h78a, 12'h669, 12'h669, 12'h569, 12'h569, 12'h67a, 12'h78a, 12'h88b, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcbd, 12'hcbd, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'hbbd, 12'haac, 12'h99b, 12'h88a, 12'h88a, 12'h889, 12'h889, 
12'h98a, 12'ha9b, 12'haac, 12'hbbc, 12'hcbc, 12'hccd, 12'hccd, 12'hbbb, 12'h779, 12'h557, 12'h346, 12'h446, 12'h557, 12'h678, 12'h668, 12'h567, 12'h567, 12'h667, 12'h668, 12'h668, 12'h668, 12'h668, 12'h679, 12'h779, 12'h88a, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heed, 12'hddd, 12'hbbb, 12'h999, 12'h777, 12'h665, 12'h554, 12'h554, 12'h444, 12'h433, 12'h322, 12'h433, 12'h544, 12'h544, 12'h434, 12'h334, 12'h325, 12'h226, 12'h226, 12'h227, 12'h337, 12'h348, 12'h458, 12'h569, 12'h67a, 12'h77b, 12'h78b, 12'h88c, 12'h89c, 12'h99d, 12'h99d, 12'h99d, 12'h9ad, 12'haad, 12'haad, 12'haad, 12'hbad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hcbe, 12'hcbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hccd, 12'hbbd, 
12'h9ac, 12'h89b, 12'h67a, 12'h569, 12'h569, 12'h569, 12'h669, 12'h67a, 12'h78b, 12'h89c, 12'h9ac, 12'hbbd, 12'hbce, 12'hcce, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hcbd, 12'hbbd, 12'haac, 12'haab, 12'ha9b, 12'ha9b, 12'haab, 12'haab, 
12'hbbc, 12'hbbc, 12'hccd, 12'hdcd, 12'hdde, 12'hdde, 12'hdde, 12'hbbc, 12'h88a, 12'h667, 12'h446, 12'h456, 12'h567, 12'h678, 12'h678, 12'h567, 12'h557, 12'h567, 12'h567, 12'h668, 12'h668, 12'h668, 12'h679, 12'h779, 12'h88a, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hddd, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccb, 12'haa9, 12'h887, 12'h666, 12'h554, 12'h554, 12'h544, 12'h433, 12'h322, 12'h433, 12'h544, 12'h544, 12'h433, 12'h324, 12'h325, 12'h226, 12'h337, 12'h337, 12'h347, 12'h458, 12'h569, 12'h66a, 12'h77b, 12'h88b, 12'h89c, 12'h99c, 12'h99d, 12'h9ad, 12'haad, 12'haae, 12'haae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hbbd, 12'haac, 
12'h99b, 12'h88a, 12'h669, 12'h559, 12'h569, 12'h569, 12'h67a, 12'h77a, 12'h88b, 12'h99c, 12'haad, 12'hbbd, 12'hbce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hcbd, 12'hbbd, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hcbd, 12'hccd, 
12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hdde, 12'hdde, 12'hccd, 12'h99a, 12'h668, 12'h557, 12'h557, 12'h667, 12'h778, 12'h678, 12'h567, 12'h557, 12'h557, 12'h567, 12'h668, 12'h668, 12'h668, 12'h779, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'hfee, 12'hffe, 12'hffe, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccb, 12'haa9, 12'h888, 12'h776, 12'h555, 12'h554, 12'h544, 12'h433, 12'h323, 12'h433, 12'h444, 12'h444, 12'h333, 12'h323, 12'h335, 12'h336, 12'h337, 12'h447, 12'h458, 12'h569, 12'h67a, 12'h77b, 12'h88b, 12'h99c, 12'h9ad, 12'haad, 12'habe, 12'hbbe, 12'hbbe, 12'hbbf, 12'hbcf, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcce, 12'hbbd, 12'haac, 
12'h88b, 12'h77a, 12'h569, 12'h458, 12'h559, 12'h569, 12'h67a, 12'h78b, 12'h89c, 12'h9ac, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hdde, 12'hdde, 12'hccd, 12'h99a, 12'h678, 12'h557, 12'h557, 12'h667, 12'h678, 12'h678, 12'h567, 12'h557, 12'h557, 12'h557, 12'h568, 12'h668, 12'h668, 12'h678, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hffe, 12'hffe, 12'hfee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccb, 12'haaa, 12'h888, 12'h776, 12'h655, 12'h555, 12'h554, 12'h444, 12'h333, 12'h433, 12'h434, 12'h433, 12'h333, 12'h324, 12'h335, 12'h336, 12'h347, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h89c, 12'h9ad, 12'haad, 12'habe, 12'hbbe, 12'hbbe, 12'hbcf, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcce, 12'hbbd, 12'h99b, 
12'h77a, 12'h669, 12'h458, 12'h448, 12'h459, 12'h569, 12'h67a, 12'h88b, 12'h99c, 12'haad, 12'habd, 12'hbbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 
12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hccd, 12'h99a, 12'h778, 12'h557, 12'h557, 12'h667, 12'h668, 12'h668, 12'h668, 12'h567, 12'h557, 12'h557, 12'h568, 12'h668, 12'h668, 12'h668, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hddd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddc, 12'hcbb, 12'haaa, 12'h988, 12'h776, 12'h655, 12'h655, 12'h544, 12'h444, 12'h433, 12'h333, 12'h333, 12'h333, 12'h333, 12'h334, 12'h325, 12'h226, 12'h337, 12'h347, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h89c, 12'h9ad, 12'haad, 12'haae, 12'hbbe, 12'hbbe, 12'hbbf, 12'hccf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcce, 12'hbac, 12'h88b, 
12'h669, 12'h558, 12'h348, 12'h348, 12'h458, 12'h559, 12'h67a, 12'h88b, 12'h99c, 12'haad, 12'hbbd, 12'hbce, 12'hcce, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hbbd, 12'h99b, 12'h779, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h557, 12'h557, 12'h568, 12'h668, 12'h668, 12'h668, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hbcc, 12'hddd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h998, 12'h777, 12'h665, 12'h655, 12'h544, 12'h444, 12'h433, 12'h333, 12'h323, 12'h333, 12'h434, 12'h434, 12'h325, 12'h226, 12'h337, 12'h347, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99c, 12'h9ad, 12'haad, 12'haae, 12'hbbe, 12'hbbe, 12'hbbf, 12'hbcf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hdde, 12'hcbd, 12'haac, 12'h88a, 
12'h558, 12'h448, 12'h337, 12'h348, 12'h458, 12'h559, 12'h77a, 12'h89b, 12'h9ac, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hcce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hbbd, 12'haab, 12'h88a, 12'h779, 12'h678, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h668, 12'h557, 12'h558, 12'h668, 12'h668, 12'h678, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'hbaa, 12'h999, 12'h888, 12'h666, 12'h655, 12'h544, 12'h444, 12'h434, 12'h333, 12'h222, 12'h323, 12'h434, 12'h445, 12'h335, 12'h226, 12'h337, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99c, 12'h9ad, 12'haad, 12'haad, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hdde, 12'hdce, 12'hbbd, 12'h99b, 12'h779, 
12'h558, 12'h448, 12'h337, 12'h348, 12'h458, 12'h569, 12'h77a, 12'h89b, 12'h9ac, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hccd, 12'haab, 12'h99a, 12'h88a, 12'h779, 12'h778, 12'h668, 12'h668, 12'h668, 12'h668, 12'h567, 12'h557, 12'h667, 12'h668, 12'h668, 12'h778, 12'h889, 12'h99a, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'hedd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h988, 12'h777, 12'h666, 12'h545, 12'h444, 12'h444, 12'h433, 12'h222, 12'h323, 12'h434, 12'h445, 12'h336, 12'h226, 12'h337, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99c, 12'h99d, 12'haad, 12'haad, 12'haae, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hdef, 12'hdef, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hdde, 12'hccd, 12'hbac, 12'h98a, 12'h669, 
12'h558, 12'h447, 12'h337, 12'h348, 12'h558, 12'h569, 12'h77a, 12'h89c, 12'h9ac, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hbbc, 12'haab, 12'h99a, 12'h88a, 12'h779, 12'h558, 12'h557, 12'h658, 12'h668, 12'h557, 12'h557, 12'h557, 12'h668, 12'h668, 12'h778, 12'h889, 12'h99a, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbba, 12'h999, 12'h888, 12'h766, 12'h555, 12'h444, 12'h444, 12'h434, 12'h323, 12'h323, 12'h434, 12'h445, 12'h336, 12'h336, 12'h337, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99c, 12'h9ad, 12'haad, 12'haad, 12'haae, 12'habe, 12'hbbe, 12'hbbe, 12'hbbf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'heef, 12'hedf, 12'hdce, 12'hbbc, 12'ha9b, 12'h879, 12'h668, 
12'h558, 12'h447, 12'h347, 12'h448, 12'h559, 12'h669, 12'h78a, 12'h89c, 12'h9ac, 12'habd, 12'hbbe, 12'hcce, 12'hccf, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hbbc, 12'haab, 12'h99a, 12'h879, 12'h668, 12'h558, 12'h668, 12'h668, 12'h557, 12'h547, 12'h557, 12'h668, 12'h778, 12'h889, 12'h989, 12'h99a, 12'haab, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h767, 12'h555, 12'h545, 12'h545, 12'h444, 12'h333, 12'h323, 12'h434, 12'h435, 12'h325, 12'h226, 12'h337, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h99c, 12'h9ad, 12'haad, 12'haae, 12'haae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hede, 12'hedf, 12'hfef, 12'hedf, 12'hccd, 12'hbac, 12'h98a, 12'h769, 12'h558, 
12'h558, 12'h558, 12'h448, 12'h458, 12'h569, 12'h67a, 12'h78b, 12'h89c, 12'h9ac, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'hccd, 12'hbbc, 12'haab, 12'h88a, 12'h779, 12'h668, 12'h779, 12'h779, 12'h658, 12'h557, 12'h667, 12'h778, 12'h779, 12'h889, 12'h99a, 12'haab, 12'hbbb, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heed, 12'hddd, 12'hddc, 12'hcbb, 12'haaa, 12'h888, 12'h777, 12'h555, 12'h545, 12'h545, 12'h445, 12'h434, 12'h334, 12'h434, 12'h435, 12'h325, 12'h226, 12'h337, 12'h437, 12'h558, 12'h669, 12'h77a, 12'h88b, 12'h89c, 12'h99d, 12'h9ad, 12'haad, 12'haae, 12'habe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbf, 12'hccf, 12'hccf, 12'hccf, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hedf, 12'heef, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'hedf, 12'heef, 12'hfef, 12'hede, 12'hcbd, 12'ha9b, 12'h879, 12'h658, 12'h547, 
12'h558, 12'h558, 12'h448, 12'h458, 12'h569, 12'h67a, 12'h77a, 12'h88b, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 
12'hddf, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hbac, 12'h99b, 12'h88a, 12'h879, 12'h88a, 12'h879, 12'h668, 12'h557, 12'h668, 12'h778, 12'h889, 12'h99a, 12'haaa, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hdcc, 12'hbbb, 12'haaa, 12'h888, 12'h766, 12'h555, 12'h544, 12'h545, 12'h545, 12'h434, 12'h434, 12'h434, 12'h334, 12'h225, 12'h226, 12'h226, 12'h337, 12'h448, 12'h569, 12'h67a, 12'h77b, 12'h88c, 12'h99c, 12'h99d, 12'haad, 12'haae, 12'haae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcbe, 12'hccf, 12'hccf, 12'hdcf, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'hede, 12'hbbc, 12'h98a, 12'h769, 12'h657, 12'h547, 
12'h558, 12'h558, 12'h548, 12'h558, 12'h669, 12'h66a, 12'h77a, 12'h88b, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hbbc, 12'ha9b, 12'h99b, 12'haab, 12'h99b, 12'h879, 12'h668, 12'h778, 12'h889, 12'h99a, 12'haab, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h888, 12'h666, 12'h555, 12'h444, 12'h545, 12'h545, 12'h445, 12'h434, 12'h434, 12'h334, 12'h225, 12'h226, 12'h226, 12'h337, 12'h448, 12'h559, 12'h66a, 12'h77a, 12'h88b, 12'h89c, 12'h99d, 12'h99d, 12'haad, 12'haae, 12'hbae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hede, 12'hede, 12'hdcd, 12'hbab, 12'h879, 12'h768, 12'h547, 12'h547, 
12'h557, 12'h558, 12'h448, 12'h448, 12'h559, 12'h669, 12'h67a, 12'h77b, 12'h88b, 12'h9ac, 12'habd, 12'hbbe, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdce, 12'hccd, 12'hbbd, 12'hbbc, 12'hbbd, 12'hbbc, 12'h99a, 12'h779, 12'h889, 12'ha9a, 12'haab, 12'hbbc, 12'hccc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'ha99, 12'h888, 12'h767, 12'h655, 12'h545, 12'h545, 12'h545, 12'h445, 12'h434, 12'h434, 12'h434, 12'h335, 12'h336, 12'h337, 12'h337, 12'h448, 12'h559, 12'h669, 12'h77a, 12'h78b, 12'h88c, 12'h99c, 12'h99d, 12'haad, 12'haae, 12'haae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hede, 12'hdcd, 12'hcbc, 12'ha8a, 12'h768, 12'h657, 12'h547, 12'h547, 
12'h547, 12'h547, 12'h447, 12'h448, 12'h448, 12'h558, 12'h559, 12'h66a, 12'h77b, 12'h89c, 12'haad, 12'hbbd, 12'hbce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hddf, 12'hddf, 12'hedf, 12'hddf, 12'hdde, 12'hdce, 12'hccd, 12'hccd, 12'hccd, 12'hcbd, 12'h99b, 12'h88a, 12'h99a, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h988, 12'h777, 12'h666, 12'h555, 12'h545, 12'h545, 12'h445, 12'h445, 12'h434, 12'h434, 12'h335, 12'h336, 12'h337, 12'h337, 12'h448, 12'h559, 12'h669, 12'h67a, 12'h77b, 12'h88c, 12'h99c, 12'h99d, 12'h9ad, 12'haad, 12'haae, 12'hbae, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hede, 12'hcbc, 12'hb9b, 12'h979, 12'h757, 12'h647, 12'h547, 12'h547, 
12'h547, 12'h547, 12'h447, 12'h447, 12'h448, 12'h448, 12'h448, 12'h559, 12'h66a, 12'h78b, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'heef, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdce, 12'hdce, 12'hdce, 12'hccd, 12'ha9b, 12'h88a, 12'h99a, 12'hbbc, 12'hccd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h777, 12'h656, 12'h545, 12'h445, 12'h434, 12'h434, 12'h434, 12'h334, 12'h325, 12'h326, 12'h327, 12'h337, 12'h337, 12'h448, 12'h559, 12'h66a, 12'h77b, 12'h88b, 12'h88c, 12'h99c, 12'h99d, 12'haad, 12'haae, 12'haae, 12'hbae, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hede, 12'hdcd, 12'hbab, 12'h989, 12'h868, 12'h647, 12'h647, 12'h647, 12'h547, 
12'h437, 12'h437, 12'h437, 12'h337, 12'h227, 12'h227, 12'h238, 12'h348, 12'h559, 12'h66a, 12'h88b, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hcdf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'heef, 
12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hddf, 12'hedf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdce, 12'hccd, 12'ha9b, 12'h98a, 12'haab, 12'hccd, 12'hddd, 12'hede, 12'heee, 12'heee, 12'hfef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hcbb, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h667, 12'h555, 12'h445, 12'h434, 12'h434, 12'h334, 12'h324, 12'h325, 12'h326, 12'h226, 12'h226, 12'h327, 12'h448, 12'h459, 12'h559, 12'h66a, 12'h77b, 12'h88c, 12'h88c, 12'h99d, 12'h99d, 12'haad, 12'haae, 12'hbae, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hede, 12'hede, 12'hcbc, 12'ha9a, 12'h868, 12'h657, 12'h546, 12'h546, 12'h647, 12'h547, 
12'h436, 12'h436, 12'h336, 12'h336, 12'h226, 12'h227, 12'h227, 12'h338, 12'h448, 12'h559, 12'h77a, 12'h88b, 12'h99c, 12'haad, 12'hbbd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 
12'hdef, 12'heef, 12'hdef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'heef, 12'heef, 12'hede, 12'hede, 12'hede, 12'hdde, 12'hccd, 12'hbbc, 12'ha9b, 12'ha9a, 12'hbbc, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hcbb, 12'hbbb, 12'haaa, 12'h888, 12'h777, 12'h655, 12'h544, 12'h434, 12'h434, 12'h423, 12'h424, 12'h325, 12'h326, 12'h326, 12'h326, 12'h327, 12'h437, 12'h448, 12'h559, 12'h66a, 12'h77b, 12'h77b, 12'h88c, 12'h98c, 12'h99d, 12'h99d, 12'haad, 12'haae, 12'hbae, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddd, 12'hccc, 12'hbab, 12'h989, 12'h767, 12'h646, 12'h535, 12'h546, 12'h546, 12'h546, 
12'h546, 12'h446, 12'h435, 12'h436, 12'h336, 12'h336, 12'h336, 12'h437, 12'h447, 12'h558, 12'h669, 12'h77a, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hcdf, 12'hcce, 12'hcce, 12'hcce, 12'hbce, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 
12'hddf, 12'hdef, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heef, 12'heef, 12'heef, 12'heee, 12'hede, 12'heee, 12'heef, 12'hdde, 12'hcbc, 12'hbab, 12'haaa, 12'hbab, 12'hccc, 12'heed, 12'heee, 12'heee, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hedd, 12'hddd, 12'hccc, 12'hcbb, 12'hbaa, 12'h999, 12'h877, 12'h665, 12'h544, 12'h533, 12'h433, 12'h423, 12'h423, 12'h424, 12'h426, 12'h426, 12'h436, 12'h437, 12'h537, 12'h548, 12'h559, 12'h669, 12'h76a, 12'h77b, 12'h87b, 12'h88c, 12'h99c, 12'h99d, 12'ha9d, 12'haad, 12'haad, 12'hbae, 12'hbbe, 12'hbbe, 12'hcce, 12'hccf, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcde, 12'hccd, 12'haab, 12'h999, 12'h878, 12'h656, 12'h545, 12'h434, 12'h445, 12'h545, 12'h545, 
12'h545, 12'h445, 12'h435, 12'h435, 12'h435, 12'h446, 12'h446, 12'h446, 12'h446, 12'h446, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcdf, 12'hccf, 12'hcce, 12'hcce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 
12'hddf, 12'hddf, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hcbc, 12'hbab, 12'hbab, 12'hbbc, 12'hdcd, 12'heee, 12'heee, 12'hfee, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'hddd, 12'hdcc, 12'hccb, 12'hbaa, 12'h999, 12'h877, 12'h765, 12'h654, 12'h533, 12'h533, 12'h533, 12'h533, 12'h534, 12'h425, 12'h426, 12'h436, 12'h436, 12'h537, 12'h547, 12'h548, 12'h659, 12'h66a, 12'h76a, 12'h77b, 12'h88b, 12'h88c, 12'h99c, 12'h99d, 12'haad, 12'haad, 12'haad, 12'hbad, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hbbc, 12'ha9a, 12'h888, 12'h767, 12'h656, 12'h445, 12'h434, 12'h434, 12'h545, 12'h445, 
12'h445, 12'h435, 12'h435, 12'h435, 12'h445, 12'h446, 12'h446, 12'h446, 12'h446, 12'h336, 12'h446, 12'h557, 12'h668, 12'h889, 12'h99a, 12'haab, 12'hbbc, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcbd, 12'hbbd, 12'hbbd, 12'haad, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hddf, 12'hdef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcdf, 12'hccf, 12'hcce, 12'hbce, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hccf, 12'hccf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 
12'hddf, 12'hddf, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heee, 12'hede, 12'hdcd, 12'hcbc, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'hfee, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'hddd, 12'hdcc, 12'hcbb, 12'hbaa, 12'h998, 12'h776, 12'h655, 12'h544, 12'h543, 12'h543, 12'h544, 12'h544, 12'h535, 12'h425, 12'h425, 12'h425, 12'h436, 12'h436, 12'h437, 12'h548, 12'h558, 12'h659, 12'h66a, 12'h77a, 12'h77b, 12'h88c, 12'h99c, 12'h99d, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbe, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hbcd, 12'hbcd, 12'haab, 12'h989, 12'h777, 12'h656, 12'h545, 12'h434, 12'h334, 12'h434, 12'h434, 12'h434, 
12'h434, 12'h334, 12'h335, 12'h435, 12'h445, 12'h446, 12'h446, 12'h436, 12'h336, 12'h225, 12'h336, 12'h447, 12'h558, 12'h779, 12'h88a, 12'h99b, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'ha9c, 12'h99b, 12'h99b, 12'haac, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcdf, 12'hcdf, 12'hcce, 12'hcce, 12'hbbe, 12'hbbd, 12'habd, 12'hbbd, 12'hbbe, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 
12'hdde, 12'hddf, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'hede, 12'hddd, 12'hccc, 12'hbbc, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hdcc, 12'hcbb, 12'hbaa, 12'h998, 12'h776, 12'h655, 12'h544, 12'h533, 12'h543, 12'h544, 12'h645, 12'h545, 12'h435, 12'h425, 12'h425, 12'h426, 12'h436, 12'h437, 12'h447, 12'h548, 12'h559, 12'h669, 12'h66a, 12'h77b, 12'h88b, 12'h88c, 12'h99c, 12'h99d, 12'haad, 12'haad, 12'haad, 12'hbad, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'habc, 12'h99b, 12'h778, 12'h666, 12'h545, 12'h444, 12'h433, 12'h333, 12'h434, 12'h444, 12'h434, 
12'h334, 12'h334, 12'h334, 12'h435, 12'h445, 12'h446, 12'h446, 12'h336, 12'h335, 12'h225, 12'h225, 12'h336, 12'h447, 12'h558, 12'h668, 12'h779, 12'h88a, 12'h98b, 12'h99b, 12'haac, 12'haac, 12'haac, 12'h99c, 12'h88b, 12'h87a, 12'h669, 12'h669, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hcce, 12'hcde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcce, 12'hcce, 12'hbce, 12'hbbd, 12'habd, 12'habd, 12'hbbd, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 
12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heef, 12'hede, 12'hdcd, 12'hcbc, 12'hbbb, 12'hbbb, 12'hccd, 12'hede, 12'heee, 12'hfee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hedd, 12'hddc, 12'hccb, 12'hbaa, 12'h999, 12'h877, 12'h665, 12'h544, 12'h533, 12'h543, 12'h544, 12'h544, 12'h544, 12'h434, 12'h425, 12'h425, 12'h425, 12'h436, 12'h436, 12'h437, 12'h448, 12'h558, 12'h559, 12'h66a, 12'h77a, 12'h87b, 12'h88c, 12'h99c, 12'h99d, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'habc, 12'h9ac, 12'h88a, 12'h667, 12'h554, 12'h443, 12'h333, 12'h433, 12'h333, 12'h444, 12'h444, 12'h444, 
12'h334, 12'h334, 12'h334, 12'h445, 12'h445, 12'h445, 12'h446, 12'h335, 12'h335, 12'h336, 12'h336, 12'h336, 12'h336, 12'h336, 12'h447, 12'h558, 12'h668, 12'h779, 12'h88a, 12'h99b, 12'h99b, 12'h99c, 12'h99b, 12'h88b, 12'h76a, 12'h549, 12'h448, 12'h659, 12'h769, 12'h88a, 12'h99b, 12'hbbc, 12'hccd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcce, 12'hcce, 12'hbbd, 12'habd, 12'haad, 12'haad, 12'habd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hccc, 12'hbbc, 12'hbbb, 12'hcbc, 12'hdcd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hbbb, 12'ha99, 12'h887, 12'h766, 12'h654, 12'h533, 12'h433, 12'h543, 12'h544, 12'h534, 12'h434, 12'h434, 12'h434, 12'h435, 12'h435, 12'h436, 12'h436, 12'h447, 12'h448, 12'h559, 12'h669, 12'h66a, 12'h77b, 12'h88b, 12'h98c, 12'h99c, 12'ha9d, 12'haad, 12'haad, 12'hbad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'haac, 12'h89b, 12'h779, 12'h556, 12'h444, 12'h333, 12'h333, 12'h343, 12'h444, 12'h444, 12'h444, 12'h444, 
12'h344, 12'h344, 12'h344, 12'h445, 12'h445, 12'h445, 12'h445, 12'h335, 12'h336, 12'h446, 12'h446, 12'h336, 12'h336, 12'h336, 12'h337, 12'h447, 12'h558, 12'h769, 12'h88a, 12'h99b, 12'haac, 12'haac, 12'haac, 12'h99c, 12'h98b, 12'h77a, 12'h669, 12'h669, 12'h669, 12'h779, 12'h99b, 12'haac, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hdef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcde, 12'hcce, 12'hbbd, 12'habd, 12'haac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'hede, 12'hddd, 12'hcbc, 12'hbbb, 12'hbbc, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'hddd, 12'hddc, 12'hcbb, 12'haaa, 12'h988, 12'h776, 12'h655, 12'h533, 12'h432, 12'h533, 12'h533, 12'h433, 12'h433, 12'h434, 12'h434, 12'h435, 12'h435, 12'h436, 12'h436, 12'h447, 12'h447, 12'h458, 12'h559, 12'h66a, 12'h77b, 12'h88b, 12'h88c, 12'h99c, 12'h99c, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbad, 12'haad, 12'haac, 12'haac, 12'habd, 12'hbbd, 12'hbbd, 12'habd, 12'h9ac, 12'h78a, 12'h668, 12'h455, 12'h344, 12'h343, 12'h344, 12'h444, 12'h454, 12'h455, 12'h455, 12'h455, 
12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h445, 12'h345, 12'h335, 12'h446, 12'h446, 12'h447, 12'h447, 12'h446, 12'h336, 12'h336, 12'h447, 12'h558, 12'h779, 12'h88b, 12'haac, 12'hbbd, 12'hcbd, 12'hcce, 12'hbbd, 12'hbbd, 12'haac, 12'h99b, 12'h779, 12'h668, 12'h779, 12'h88a, 12'ha9b, 12'hbbc, 12'hccd, 12'hdde, 12'hdef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hcce, 12'hbcd, 12'habd, 12'haac, 12'h99c, 12'h99b, 12'h99c, 12'haac, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdde, 12'hdcd, 12'hcbc, 12'hbbb, 12'hcbc, 12'hccc, 12'hede, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hbba, 12'h999, 12'h877, 12'h655, 12'h533, 12'h421, 12'h432, 12'h433, 12'h433, 12'h433, 12'h434, 12'h444, 12'h445, 12'h445, 12'h445, 12'h336, 12'h346, 12'h447, 12'h448, 12'h559, 12'h669, 12'h77a, 12'h77b, 12'h88b, 12'h88c, 12'h99c, 12'h99c, 12'haad, 12'haad, 12'haac, 12'ha9c, 12'ha9c, 12'h99c, 12'ha9c, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'habd, 12'habd, 12'haac, 12'h99b, 12'h78a, 12'h568, 12'h456, 12'h344, 12'h344, 12'h344, 12'h444, 12'h454, 12'h455, 12'h455, 12'h455, 
12'h445, 12'h445, 12'h345, 12'h335, 12'h345, 12'h345, 12'h345, 12'h346, 12'h446, 12'h446, 12'h447, 12'h447, 12'h557, 12'h557, 12'h558, 12'h668, 12'h679, 12'h88a, 12'h99b, 12'haac, 12'hcbd, 12'hcce, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hbbd, 12'haab, 12'h99b, 12'h99b, 12'haab, 12'hbac, 12'hbbd, 12'hcce, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hddf, 12'hddf, 12'hddf, 12'hdef, 12'hddf, 12'hdde, 12'hcce, 12'hbbd, 12'haac, 12'h9ac, 12'h99b, 12'h99b, 12'h99c, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'hede, 12'hddd, 12'hccd, 12'hcbc, 12'hcbc, 12'hccc, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hbbb, 12'ha99, 12'h877, 12'h665, 12'h533, 12'h421, 12'h433, 12'h533, 12'h443, 12'h443, 12'h443, 12'h444, 12'h444, 12'h445, 12'h445, 12'h345, 12'h346, 12'h347, 12'h447, 12'h458, 12'h569, 12'h66a, 12'h77a, 12'h78b, 12'h88b, 12'h88b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h98c, 12'h98b, 12'h98b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haac, 12'haac, 12'h99b, 12'h78a, 12'h668, 12'h556, 12'h445, 12'h344, 12'h344, 12'h344, 12'h334, 12'h344, 12'h345, 12'h345, 
12'h345, 12'h335, 12'h334, 12'h224, 12'h235, 12'h235, 12'h335, 12'h446, 12'h446, 12'h346, 12'h446, 12'h557, 12'h668, 12'h779, 12'h779, 12'h88a, 12'h88a, 12'h99b, 12'haac, 12'hbbc, 12'hccd, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hdef, 12'hddf, 12'hdde, 12'hccd, 12'hbbd, 12'haac, 12'h99b, 12'h88b, 12'h89b, 12'h99b, 12'haac, 12'haad, 12'hbbd, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hccd, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hede, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hbbb, 12'ha99, 12'h887, 12'h766, 12'h543, 12'h422, 12'h533, 12'h543, 12'h543, 12'h443, 12'h443, 12'h444, 12'h444, 12'h445, 12'h445, 12'h345, 12'h346, 12'h346, 12'h347, 12'h448, 12'h559, 12'h669, 12'h66a, 12'h77a, 12'h77b, 12'h87b, 12'h88b, 12'h98b, 12'h98b, 12'h88b, 12'h87b, 12'h87a, 12'h87a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'h99b, 12'h78a, 12'h679, 12'h567, 12'h456, 12'h445, 12'h335, 12'h234, 12'h124, 12'h234, 12'h235, 12'h235, 
12'h235, 12'h235, 12'h224, 12'h124, 12'h225, 12'h235, 12'h346, 12'h446, 12'h447, 12'h446, 12'h457, 12'h668, 12'h779, 12'h88a, 12'h99a, 12'h9ab, 12'haab, 12'haac, 12'hbbc, 12'hbbd, 12'hccd, 12'hcde, 12'hdde, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hede, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hcde, 12'hccd, 12'habc, 12'h99b, 12'h88b, 12'h88a, 12'h88a, 12'h88b, 12'h99c, 12'haac, 12'hbbd, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'heef, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hede, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hdcc, 12'hcbb, 12'haa9, 12'h988, 12'h766, 12'h544, 12'h432, 12'h533, 12'h544, 12'h543, 12'h442, 12'h443, 12'h453, 12'h444, 12'h444, 12'h445, 12'h345, 12'h335, 12'h346, 12'h347, 12'h447, 12'h458, 12'h569, 12'h669, 12'h66a, 12'h77a, 12'h77a, 12'h77b, 12'h88b, 12'h88b, 12'h87a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h87a, 12'h77a, 12'h77a, 12'h87a, 12'h88b, 12'h89b, 12'h99c, 12'h9ac, 12'h89b, 12'h88b, 12'h779, 12'h668, 12'h567, 12'h556, 12'h446, 12'h345, 12'h235, 12'h235, 12'h335, 12'h346, 
12'h346, 12'h346, 12'h336, 12'h336, 12'h346, 12'h446, 12'h557, 12'h668, 12'h778, 12'h779, 12'h889, 12'h99a, 12'h9ab, 12'haac, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hbcd, 12'hccd, 12'hccd, 12'hcde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hcde, 12'hccd, 12'haac, 12'h99b, 12'h88a, 12'h77a, 12'h77a, 12'h88a, 12'h99b, 12'haac, 12'hbbd, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdce, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'hdcd, 12'hddd, 12'heee, 12'hfee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hddd, 12'hddc, 12'hccb, 12'hbaa, 12'h998, 12'h776, 12'h544, 12'h422, 12'h533, 12'h543, 12'h543, 12'h442, 12'h442, 12'h453, 12'h444, 12'h444, 12'h345, 12'h345, 12'h235, 12'h236, 12'h336, 12'h447, 12'h558, 12'h569, 12'h669, 12'h66a, 12'h66a, 12'h77a, 12'h77a, 12'h87b, 12'h87b, 12'h77a, 12'h77a, 12'h77a, 12'h76a, 12'h77a, 12'h77a, 12'h779, 12'h769, 12'h779, 12'h77a, 12'h78a, 12'h88b, 12'h99b, 12'h89b, 12'h88b, 12'h78a, 12'h779, 12'h779, 12'h668, 12'h668, 12'h557, 12'h457, 12'h457, 12'h457, 12'h557, 
12'h568, 12'h568, 12'h568, 12'h568, 12'h668, 12'h678, 12'h779, 12'h88a, 12'h99a, 12'haab, 12'haac, 12'hbbc, 12'hbcd, 12'hccd, 12'hccd, 12'hcdd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heef, 12'hfef, 12'hfef, 12'hfef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'hdef, 12'hdee, 12'hdde, 12'hcce, 12'hbbd, 12'haab, 12'h88a, 12'h779, 12'h669, 12'h669, 12'h88a, 12'h99c, 12'haad, 12'hbbd, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hddd, 12'hccc, 12'hccd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hedd, 12'hddd, 12'hccc, 12'hbba, 12'ha99, 12'h877, 12'h654, 12'h422, 12'h533, 12'h433, 12'h442, 12'h442, 12'h442, 12'h453, 12'h444, 12'h444, 12'h444, 12'h345, 12'h235, 12'h346, 12'h347, 12'h457, 12'h558, 12'h569, 12'h669, 12'h67a, 12'h77a, 12'h77a, 12'h77a, 12'h87a, 12'h87a, 12'h77a, 12'h77a, 12'h769, 12'h769, 12'h769, 12'h769, 12'h669, 12'h669, 12'h669, 12'h669, 12'h779, 12'h78a, 12'h88b, 12'h88b, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h779, 12'h779, 12'h679, 12'h679, 12'h779, 12'h779, 
12'h779, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h89a, 12'h99b, 12'haac, 12'hbbc, 12'hbbd, 12'hccd, 12'hccd, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddd, 12'hcdd, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'heef, 12'hdde, 12'hccd, 12'habc, 12'h99b, 12'h77a, 12'h569, 12'h558, 12'h669, 12'h88a, 12'h99c, 12'haac, 12'haad, 12'hbad, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdcf, 12'hddf, 12'hdce, 12'hdde, 12'hdde, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddd, 12'hdcd, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'hedd, 12'hddc, 12'hcbb, 12'haa9, 12'h888, 12'h655, 12'h422, 12'h432, 12'h432, 12'h432, 12'h442, 12'h442, 12'h443, 12'h443, 12'h444, 12'h344, 12'h345, 12'h345, 12'h346, 12'h447, 12'h458, 12'h569, 12'h679, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h87a, 12'h88a, 12'h88a, 12'h87a, 12'h77a, 12'h769, 12'h669, 12'h669, 12'h669, 12'h668, 12'h658, 12'h558, 12'h558, 12'h669, 12'h779, 12'h78a, 12'h78a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h88b, 12'h88b, 12'h99b, 12'h99b, 
12'h99b, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hccd, 12'hccd, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heee, 12'hede, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'heee, 12'heef, 12'hdde, 12'hcdd, 12'hbbd, 12'h9ab, 12'h88a, 12'h669, 12'h458, 12'h559, 12'h669, 12'h87b, 12'h99b, 12'h99c, 12'haad, 12'haad, 12'hbbd, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccf, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddd, 12'hddd, 12'hede, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'heee, 12'hddd, 12'hccc, 12'hbaa, 12'h988, 12'h765, 12'h432, 12'h432, 12'h432, 12'h431, 12'h441, 12'h442, 12'h443, 12'h443, 12'h444, 12'h344, 12'h345, 12'h345, 12'h446, 12'h457, 12'h568, 12'h679, 12'h78a, 12'h88a, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h88a, 12'h87a, 12'h77a, 12'h669, 12'h658, 12'h658, 12'h658, 12'h558, 12'h558, 12'h558, 12'h558, 12'h568, 12'h669, 12'h779, 12'h78a, 12'h78a, 12'h88a, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 
12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'heee, 12'hdde, 12'hcdd, 12'hbcd, 12'haab, 12'h88a, 12'h679, 12'h558, 12'h558, 12'h559, 12'h66a, 12'h77b, 12'h88b, 12'h99c, 12'ha9c, 12'haad, 12'hbbd, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'hedd, 12'hdcc, 12'hbbb, 12'ha99, 12'h766, 12'h543, 12'h533, 12'h432, 12'h432, 12'h442, 12'h442, 12'h443, 12'h444, 12'h444, 12'h345, 12'h345, 12'h446, 12'h457, 12'h567, 12'h678, 12'h78a, 12'h88a, 12'h89b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h88b, 12'h88a, 12'h77a, 12'h769, 12'h658, 12'h547, 12'h547, 12'h547, 12'h557, 12'h557, 12'h558, 12'h558, 12'h568, 12'h668, 12'h779, 12'h779, 12'h789, 12'h88a, 12'h99b, 12'h99c, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbad, 12'hbbd, 
12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hcdd, 12'hccd, 12'habc, 12'h99b, 12'h77a, 12'h559, 12'h558, 12'h448, 12'h559, 12'h66a, 12'h77a, 12'h88b, 12'h99c, 12'haac, 12'hbad, 12'hbbd, 12'hbbe, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'hddd, 12'hcbb, 12'haa9, 12'h876, 12'h544, 12'h543, 12'h533, 12'h432, 12'h442, 12'h442, 12'h443, 12'h444, 12'h444, 12'h445, 12'h345, 12'h446, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h99b, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'h99b, 12'h88b, 12'h88a, 12'h779, 12'h669, 12'h547, 12'h436, 12'h436, 12'h436, 12'h447, 12'h557, 12'h557, 12'h557, 12'h567, 12'h668, 12'h678, 12'h779, 12'h789, 12'h78a, 12'h88b, 12'h99b, 12'ha9c, 12'haad, 12'hbad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 
12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hccd, 12'hbbd, 12'haac, 12'h88a, 12'h669, 12'h558, 12'h338, 12'h448, 12'h559, 12'h66a, 12'h77a, 12'h88b, 12'h99c, 12'haac, 12'haad, 12'hbbd, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hddd, 12'hccc, 12'hbaa, 12'h877, 12'h644, 12'h544, 12'h543, 12'h443, 12'h433, 12'h433, 12'h433, 12'h434, 12'h334, 12'h335, 12'h345, 12'h456, 12'h668, 12'h779, 12'h88a, 12'h9ab, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'haac, 12'haac, 12'h99b, 12'h88a, 12'h669, 12'h558, 12'h447, 12'h436, 12'h436, 12'h436, 12'h446, 12'h446, 12'h456, 12'h446, 12'h456, 12'h567, 12'h668, 12'h678, 12'h778, 12'h789, 12'h88a, 12'h88b, 12'h99c, 12'haac, 12'haad, 12'haad, 12'hbad, 12'hbbd, 12'hbbd, 
12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'hfef, 12'hfef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hccd, 12'hbbc, 12'h99b, 12'h669, 12'h558, 12'h448, 12'h448, 12'h559, 12'h66a, 12'h66a, 12'h66a, 12'h87b, 12'h98c, 12'h99c, 12'haad, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'hfee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hedd, 12'hdcc, 12'hbba, 12'h887, 12'h544, 12'h543, 12'h543, 12'h543, 12'h433, 12'h433, 12'h333, 12'h333, 12'h334, 12'h335, 12'h346, 12'h557, 12'h678, 12'h88a, 12'h99b, 12'hbbc, 12'hbcd, 12'hccd, 12'hcce, 12'hccd, 12'hbbd, 12'hbbd, 12'haac, 12'h99b, 12'h668, 12'h447, 12'h436, 12'h446, 12'h436, 12'h335, 12'h335, 12'h335, 12'h335, 12'h335, 12'h345, 12'h456, 12'h567, 12'h567, 12'h677, 12'h678, 12'h77a, 12'h77a, 12'h88b, 12'h99b, 12'h99c, 12'haac, 12'haac, 12'haad, 12'hbbd, 
12'hbbd, 12'hbbd, 12'hbbd, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'hfef, 12'hfef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hbcd, 12'haab, 12'h77a, 12'h669, 12'h448, 12'h448, 12'h559, 12'h569, 12'h559, 12'h559, 12'h66a, 12'h77b, 12'h88b, 12'h99c, 12'haad, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hedd, 12'hddd, 12'hcbb, 12'h988, 12'h644, 12'h544, 12'h543, 12'h533, 12'h433, 12'h434, 12'h333, 12'h324, 12'h324, 12'h335, 12'h446, 12'h557, 12'h779, 12'h89a, 12'haac, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hbbd, 12'haac, 12'h779, 12'h557, 12'h436, 12'h436, 12'h335, 12'h335, 12'h334, 12'h334, 12'h334, 12'h234, 12'h334, 12'h345, 12'h455, 12'h456, 12'h466, 12'h567, 12'h669, 12'h679, 12'h77a, 12'h88a, 12'h88b, 12'h99b, 12'h99b, 12'h99c, 12'haac, 
12'haac, 12'haac, 12'haad, 12'hbad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hdde, 12'hccd, 12'haac, 12'h88a, 12'h779, 12'h458, 12'h348, 12'h448, 12'h448, 12'h348, 12'h348, 12'h559, 12'h66a, 12'h87b, 12'h98c, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'hfef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'hddd, 12'hcbb, 12'h988, 12'h654, 12'h544, 12'h543, 12'h543, 12'h434, 12'h434, 12'h434, 12'h434, 12'h435, 12'h435, 12'h446, 12'h657, 12'h779, 12'h89a, 12'haac, 12'hbcd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hbbc, 12'h88a, 12'h668, 12'h446, 12'h335, 12'h324, 12'h324, 12'h334, 12'h334, 12'h344, 12'h334, 12'h334, 12'h344, 12'h344, 12'h344, 12'h344, 12'h356, 12'h457, 12'h558, 12'h669, 12'h679, 12'h779, 12'h77a, 12'h88a, 12'h88a, 12'h88b, 
12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'h99c, 12'ha9c, 12'haac, 12'haac, 12'hbbd, 12'hcbe, 12'hcce, 12'hdce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hfef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hcde, 12'hbbd, 12'h99b, 12'h78a, 12'h558, 12'h348, 12'h448, 12'h348, 12'h338, 12'h338, 12'h448, 12'h559, 12'h66a, 12'h88b, 12'h99c, 12'haad, 12'hbbd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hedd, 12'hccc, 12'ha99, 12'h655, 12'h654, 12'h543, 12'h543, 12'h544, 12'h434, 12'h435, 12'h435, 12'h435, 12'h435, 12'h446, 12'h657, 12'h779, 12'h89a, 12'haac, 12'hccd, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'h99b, 12'h779, 12'h556, 12'h335, 12'h224, 12'h324, 12'h334, 12'h344, 12'h344, 12'h344, 12'h343, 12'h244, 12'h244, 12'h244, 12'h244, 12'h345, 12'h346, 12'h447, 12'h557, 12'h568, 12'h668, 12'h668, 12'h669, 12'h679, 12'h779, 
12'h77a, 12'h78a, 12'h88a, 12'h88a, 12'h88a, 12'h88b, 12'h98b, 12'h99b, 12'ha9c, 12'haad, 12'hbbd, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdce, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hbcd, 12'haac, 12'h88a, 12'h669, 12'h348, 12'h448, 12'h348, 12'h348, 12'h448, 12'h448, 12'h448, 12'h559, 12'h77a, 12'h88b, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hdcc, 12'ha99, 12'h766, 12'h765, 12'h644, 12'h534, 12'h534, 12'h435, 12'h435, 12'h435, 12'h435, 12'h435, 12'h446, 12'h557, 12'h779, 12'h88a, 12'haac, 12'hbcd, 12'hdde, 12'hddf, 12'hdef, 12'hdef, 12'hddf, 12'hdde, 12'hdde, 12'hccd, 12'haab, 12'h889, 12'h667, 12'h335, 12'h324, 12'h334, 12'h334, 12'h344, 12'h344, 12'h343, 12'h343, 12'h243, 12'h243, 12'h244, 12'h344, 12'h344, 12'h235, 12'h235, 12'h345, 12'h446, 12'h456, 12'h457, 12'h457, 12'h457, 12'h557, 
12'h558, 12'h568, 12'h668, 12'h669, 12'h669, 12'h669, 12'h77a, 12'h77a, 12'h88b, 12'h99b, 12'ha9c, 12'haad, 12'hbad, 12'hbbd, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdcf, 12'hdcf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'haac, 12'h99b, 12'h669, 12'h448, 12'h448, 12'h348, 12'h448, 12'h458, 12'h448, 12'h338, 12'h449, 12'h67a, 12'h88b, 12'h99c, 12'haad, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hdcc, 12'hbaa, 12'h877, 12'h766, 12'h644, 12'h534, 12'h534, 12'h435, 12'h435, 12'h435, 12'h435, 12'h435, 12'h436, 12'h557, 12'h669, 12'h88a, 12'haac, 12'hbbd, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hbbc, 12'h99a, 12'h767, 12'h445, 12'h334, 12'h334, 12'h344, 12'h344, 12'h343, 12'h333, 12'h233, 12'h233, 12'h243, 12'h243, 12'h354, 12'h344, 12'h133, 12'h133, 12'h234, 12'h244, 12'h245, 12'h245, 12'h245, 12'h235, 12'h345, 
12'h346, 12'h446, 12'h447, 12'h447, 12'h447, 12'h548, 12'h558, 12'h659, 12'h669, 12'h77a, 12'h87b, 12'h98b, 12'h99c, 12'ha9c, 12'haad, 12'hbad, 12'hbad, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcbe, 12'hccf, 12'hccf, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hbbd, 12'haac, 12'h99b, 12'h669, 12'h448, 12'h347, 12'h347, 12'h448, 12'h458, 12'h448, 12'h448, 12'h559, 12'h77a, 12'h88b, 12'haac, 12'habd, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hddd, 12'hbba, 12'h988, 12'h876, 12'h654, 12'h544, 12'h534, 12'h435, 12'h535, 12'h435, 12'h435, 12'h335, 12'h336, 12'h447, 12'h668, 12'h77a, 12'h99b, 12'hbbd, 12'hcce, 12'hdde, 12'hdef, 12'heef, 12'heef, 12'hddf, 12'hdde, 12'hdde, 12'hcbc, 12'haab, 12'h878, 12'h545, 12'h434, 12'h334, 12'h333, 12'h333, 12'h232, 12'h232, 12'h232, 12'h232, 12'h132, 12'h132, 12'h243, 12'h243, 12'h233, 12'h233, 12'h344, 12'h344, 12'h344, 12'h344, 12'h244, 12'h235, 12'h235, 
12'h345, 12'h346, 12'h336, 12'h336, 12'h447, 12'h447, 12'h448, 12'h548, 12'h559, 12'h659, 12'h66a, 12'h77a, 12'h87b, 12'h98b, 12'h99c, 12'ha9c, 12'ha9d, 12'haad, 12'hbad, 12'hbad, 12'hbad, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbbe, 12'hbbe, 12'hbbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hdce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hccd, 12'hbbd, 12'hbbc, 12'haac, 12'h99b, 12'h779, 12'h558, 12'h458, 12'h458, 12'h458, 12'h558, 12'h559, 12'h559, 12'h66a, 12'h88b, 12'h99c, 12'haac, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hedd, 12'hcbb, 12'ha99, 12'h877, 12'h655, 12'h544, 12'h534, 12'h535, 12'h535, 12'h435, 12'h435, 12'h325, 12'h325, 12'h436, 12'h558, 12'h779, 12'h99b, 12'hbbc, 12'hcce, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hede, 12'hdde, 12'hccd, 12'hbbc, 12'h989, 12'h656, 12'h444, 12'h334, 12'h323, 12'h222, 12'h121, 12'h121, 12'h121, 12'h122, 12'h132, 12'h132, 12'h232, 12'h232, 12'h242, 12'h242, 12'h343, 12'h344, 12'h344, 12'h344, 12'h244, 12'h234, 12'h234, 
12'h235, 12'h335, 12'h335, 12'h336, 12'h336, 12'h336, 12'h437, 12'h437, 12'h548, 12'h548, 12'h549, 12'h659, 12'h76a, 12'h77a, 12'h87b, 12'h98b, 12'h98c, 12'h99c, 12'ha9d, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haac, 12'haac, 12'haac, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbbd, 12'hcbd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbbd, 12'hbbc, 12'haac, 12'haac, 12'habc, 12'hbbc, 12'habc, 12'haab, 12'h99b, 12'h88a, 12'h78a, 12'h779, 12'h779, 12'h77a, 12'h77a, 12'h77a, 12'h78b, 12'h99b, 12'h9ac, 12'habd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heed, 12'hccc, 12'haaa, 12'h988, 12'h765, 12'h543, 12'h534, 12'h535, 12'h545, 12'h445, 12'h435, 12'h325, 12'h325, 12'h336, 12'h557, 12'h668, 12'h88a, 12'haac, 12'hbcd, 12'hcce, 12'hdde, 12'hdef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hddd, 12'hccc, 12'h99a, 12'h767, 12'h545, 12'h434, 12'h222, 12'h212, 12'h211, 12'h232, 12'h333, 12'h333, 12'h333, 12'h233, 12'h233, 12'h232, 12'h242, 12'h342, 12'h353, 12'h354, 12'h343, 12'h343, 12'h344, 12'h244, 12'h234, 
12'h334, 12'h335, 12'h335, 12'h335, 12'h326, 12'h326, 12'h327, 12'h437, 12'h437, 12'h427, 12'h428, 12'h538, 12'h549, 12'h659, 12'h65a, 12'h76a, 12'h76a, 12'h87b, 12'h98b, 12'h98c, 12'h99c, 12'h99c, 12'h99c, 12'h98c, 12'h98c, 12'h98c, 12'h98c, 12'h98b, 12'h98b, 12'h99b, 12'h99b, 12'h99b, 12'h98b, 12'h98b, 12'h99b, 12'ha9b, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haab, 12'ha9b, 12'ha9b, 12'ha9b, 12'h99b, 12'h98a, 12'h88a, 12'h99a, 12'haab, 12'habc, 12'hbbd, 12'hbbd, 12'hbbc, 12'habc, 12'haac, 12'haab, 12'haab, 12'h9ab, 12'h99b, 12'h89b, 12'h99c, 12'haac, 12'habd, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hdcc, 12'hbba, 12'h988, 12'h765, 12'h543, 12'h544, 12'h544, 12'h545, 12'h545, 12'h435, 12'h335, 12'h325, 12'h335, 12'h447, 12'h568, 12'h88a, 12'haab, 12'hbbd, 12'hccd, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hccd, 12'haab, 12'h778, 12'h656, 12'h434, 12'h323, 12'h322, 12'h322, 12'h333, 12'h444, 12'h444, 12'h444, 12'h344, 12'h334, 12'h233, 12'h342, 12'h342, 12'h453, 12'h453, 12'h453, 12'h343, 12'h344, 12'h344, 12'h344, 
12'h345, 12'h445, 12'h435, 12'h336, 12'h336, 12'h336, 12'h437, 12'h437, 12'h447, 12'h448, 12'h548, 12'h548, 12'h659, 12'h659, 12'h659, 12'h65a, 12'h76a, 12'h77a, 12'h88b, 12'h98c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h98c, 12'h98c, 12'h98b, 12'h88b, 12'h88a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h87a, 12'h88a, 12'h98b, 12'h98b, 12'h98b, 12'h98b, 12'h98a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h88a, 12'h98a, 12'h88a, 12'h88a, 12'h88a, 12'h99a, 12'haab, 12'hbbc, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbcd, 12'hbbc, 12'hbbc, 12'hbbc, 12'haac, 12'h9ac, 12'haac, 12'habd, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hcbb, 12'ha99, 12'h766, 12'h543, 12'h544, 12'h544, 12'h545, 12'h545, 12'h435, 12'h335, 12'h325, 12'h335, 12'h446, 12'h557, 12'h779, 12'h99b, 12'habc, 12'hbcd, 12'hcde, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hede, 12'hddd, 12'hbbb, 12'h989, 12'h767, 12'h545, 12'h324, 12'h323, 12'h323, 12'h334, 12'h444, 12'h445, 12'h444, 12'h344, 12'h334, 12'h333, 12'h343, 12'h342, 12'h443, 12'h443, 12'h443, 12'h343, 12'h344, 12'h344, 12'h334, 
12'h445, 12'h445, 12'h445, 12'h446, 12'h436, 12'h436, 12'h447, 12'h547, 12'h558, 12'h669, 12'h779, 12'h77a, 12'h87a, 12'h87a, 12'h77a, 12'h77a, 12'h87a, 12'h88b, 12'h99b, 12'ha9c, 12'haac, 12'haad, 12'hbad, 12'haad, 12'haac, 12'haac, 12'h99c, 12'h98b, 12'h87a, 12'h77a, 12'h669, 12'h769, 12'h77a, 12'h77a, 12'h87a, 12'h87a, 12'h87a, 12'h87a, 12'h77a, 12'h769, 12'h769, 12'h659, 12'h658, 12'h658, 12'h658, 12'h659, 12'h769, 12'h779, 12'h88a, 12'h98a, 12'h99b, 12'h99b, 12'haac, 12'hbbc, 12'hccd, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hccd, 12'hccd, 12'hccd, 12'hbcd, 12'hbbd, 12'habd, 12'hbbd, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hedd, 12'hccc, 12'haa9, 12'h766, 12'h543, 12'h544, 12'h544, 12'h544, 12'h444, 12'h434, 12'h335, 12'h334, 12'h335, 12'h346, 12'h457, 12'h678, 12'h88a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdde, 12'hcbc, 12'ha9a, 12'h878, 12'h656, 12'h434, 12'h323, 12'h213, 12'h323, 12'h334, 12'h444, 12'h445, 12'h445, 12'h345, 12'h344, 12'h343, 12'h342, 12'h342, 12'h443, 12'h443, 12'h343, 12'h333, 12'h334, 12'h334, 
12'h445, 12'h445, 12'h446, 12'h446, 12'h446, 12'h446, 12'h547, 12'h557, 12'h668, 12'h88a, 12'h99b, 12'h99b, 12'ha9b, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h99c, 12'haac, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcbd, 12'hbbd, 12'hbbd, 12'h99c, 12'h88b, 12'h77a, 12'h66a, 12'h76a, 12'h77a, 12'h88b, 12'h88b, 12'h98b, 12'h88b, 12'h87a, 12'h76a, 12'h659, 12'h548, 12'h438, 12'h427, 12'h438, 12'h538, 12'h658, 12'h769, 12'h88a, 12'h99b, 12'haac, 12'hbac, 12'hbbc, 12'hcbd, 12'hccd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcdd, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'hedd, 12'hdcc, 12'hbaa, 12'h877, 12'h654, 12'h544, 12'h544, 12'h444, 12'h444, 12'h434, 12'h334, 12'h334, 12'h235, 12'h335, 12'h446, 12'h568, 12'h789, 12'h99a, 12'haac, 12'hbcd, 12'hcde, 12'hdde, 12'hede, 12'heef, 12'heef, 12'heee, 12'hede, 12'hdcd, 12'hbbb, 12'h99a, 12'h778, 12'h556, 12'h434, 12'h323, 12'h323, 12'h324, 12'h324, 12'h334, 12'h335, 12'h335, 12'h334, 12'h333, 12'h333, 12'h443, 12'h444, 12'h444, 12'h434, 12'h333, 12'h334, 12'h334, 
12'h435, 12'h445, 12'h446, 12'h546, 12'h547, 12'h557, 12'h557, 12'h668, 12'h779, 12'h99b, 12'hbac, 12'hbbc, 12'hbbd, 12'hbbc, 12'hbac, 12'haac, 12'haac, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hbcd, 12'haac, 12'h99b, 12'h88b, 12'h77a, 12'h88b, 12'h99c, 12'haac, 12'haad, 12'haad, 12'ha9c, 12'h98b, 12'h88b, 12'h87a, 12'h76a, 12'h659, 12'h659, 12'h759, 12'h769, 12'h87a, 12'h98b, 12'ha9c, 12'hbad, 12'hcbd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcdd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heed, 12'hddd, 12'hcbb, 12'h988, 12'h766, 12'h654, 12'h543, 12'h443, 12'h443, 12'h444, 12'h334, 12'h334, 12'h334, 12'h335, 12'h346, 12'h557, 12'h779, 12'h88a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'hede, 12'hdde, 12'hccc, 12'hbab, 12'h989, 12'h778, 12'h656, 12'h545, 12'h434, 12'h324, 12'h224, 12'h224, 12'h224, 12'h335, 12'h335, 12'h444, 12'h444, 12'h545, 12'h545, 12'h445, 12'h434, 12'h334, 12'h324, 12'h325, 
12'h435, 12'h446, 12'h546, 12'h557, 12'h557, 12'h658, 12'h668, 12'h769, 12'h88a, 12'haac, 12'hcbd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hbbd, 12'hccd, 12'hccd, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hcdd, 12'hbbd, 12'haac, 12'h99b, 12'h88b, 12'h99c, 12'haad, 12'hbbe, 12'hcce, 12'hcce, 12'hbbd, 12'haad, 12'ha9c, 12'h99c, 12'h98b, 12'h87a, 12'h76a, 12'h87b, 12'h98b, 12'ha9c, 12'hbac, 12'hbbd, 12'hcce, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hcde, 12'hcdd, 12'hcdd, 12'hcdd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'hedd, 12'hccc, 12'haa9, 12'h877, 12'h665, 12'h543, 12'h443, 12'h443, 12'h443, 12'h344, 12'h334, 12'h334, 12'h335, 12'h345, 12'h456, 12'h668, 12'h789, 12'h99a, 12'hbbc, 12'hccd, 12'hdde, 12'hdde, 12'hede, 12'heef, 12'heef, 12'heee, 12'hede, 12'hddd, 12'hcbc, 12'haab, 12'h989, 12'h778, 12'h657, 12'h546, 12'h435, 12'h324, 12'h334, 12'h335, 12'h435, 12'h446, 12'h545, 12'h545, 12'h545, 12'h545, 12'h545, 12'h435, 12'h425, 12'h425, 12'h425, 
12'h436, 12'h546, 12'h547, 12'h657, 12'h658, 12'h668, 12'h768, 12'h779, 12'h98a, 12'hbbc, 12'hccd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hccd, 12'hcdd, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'heff, 12'heef, 12'heee, 12'hdee, 12'hddd, 12'hbcd, 12'haad, 12'h99c, 12'h88b, 12'h99c, 12'hbbd, 12'hcce, 12'hcce, 12'hccf, 12'hcbe, 12'hbbd, 12'haad, 12'haad, 12'ha9c, 12'h98c, 12'h98b, 12'ha9c, 12'haac, 12'hbbd, 12'hcbe, 12'hdce, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcdd, 12'hcdd, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hddc, 12'hbba, 12'h998, 12'h765, 12'h553, 12'h443, 12'h543, 12'h444, 12'h444, 12'h444, 12'h345, 12'h345, 12'h335, 12'h446, 12'h567, 12'h779, 12'h89a, 12'haab, 12'hbcd, 12'hcde, 12'hdde, 12'hede, 12'heef, 12'heee, 12'hede, 12'heee, 12'hede, 12'hdcd, 12'hcbc, 12'hbab, 12'ha9a, 12'h989, 12'h878, 12'h768, 12'h667, 12'h667, 12'h667, 12'h668, 12'h668, 12'h657, 12'h656, 12'h656, 12'h656, 12'h546, 12'h545, 12'h435, 12'h425, 12'h425, 
12'h436, 12'h546, 12'h657, 12'h657, 12'h768, 12'h779, 12'h879, 12'h889, 12'h99b, 12'hbbc, 12'hdce, 12'hdde, 12'hdde, 12'heee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heff, 12'heff, 12'heef, 12'heee, 12'hdee, 12'hcdd, 12'hbcd, 12'haad, 12'h88b, 12'h77a, 12'h88b, 12'haac, 12'hbbe, 12'hcce, 12'hcce, 12'hcbe, 12'hbbd, 12'hbad, 12'hbad, 12'hbad, 12'haad, 12'haad, 12'hbbd, 12'hcbe, 12'hcce, 12'hdcf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcdd, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hedd, 12'hccb, 12'haa9, 12'h776, 12'h654, 12'h553, 12'h554, 12'h554, 12'h444, 12'h444, 12'h445, 12'h345, 12'h345, 12'h446, 12'h557, 12'h678, 12'h88a, 12'haab, 12'hbbc, 12'hccd, 12'hdde, 12'hdde, 12'heee, 12'hede, 12'hede, 12'heee, 12'heee, 12'hede, 12'hdcd, 12'hccc, 12'hbbc, 12'hbab, 12'haab, 12'h99a, 12'h889, 12'h889, 12'h889, 12'h889, 12'h889, 12'h778, 12'h768, 12'h768, 12'h768, 12'h657, 12'h657, 12'h546, 12'h536, 12'h536, 
12'h547, 12'h547, 12'h657, 12'h658, 12'h668, 12'h779, 12'h879, 12'h88a, 12'h99b, 12'hbbc, 12'hcce, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdde, 12'hdde, 12'hdee, 12'hdee, 12'heef, 12'heff, 12'heff, 12'heff, 12'heee, 12'hdee, 12'hddd, 12'hbcd, 12'haad, 12'h88c, 12'h77b, 12'h87b, 12'h99c, 12'hbad, 12'hbbe, 12'hcce, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbad, 12'hbbd, 12'hcbe, 12'hdce, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'hfee, 12'heed, 12'hdcc, 12'hbba, 12'h887, 12'h665, 12'h554, 12'h554, 12'h544, 12'h444, 12'h444, 12'h445, 12'h445, 12'h345, 12'h446, 12'h557, 12'h668, 12'h889, 12'h9ab, 12'hbbc, 12'hccd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hccd, 12'hccd, 12'hcbd, 12'hbbc, 12'haab, 12'h99a, 12'h99a, 12'h88a, 12'h99a, 12'h98a, 12'h88a, 12'h879, 12'h779, 12'h779, 12'h769, 12'h669, 12'h668, 12'h658, 12'h558, 
12'h558, 12'h548, 12'h548, 12'h548, 12'h558, 12'h669, 12'h769, 12'h77a, 12'h99b, 12'hbbc, 12'hcce, 12'hdde, 12'hedf, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'heff, 12'heff, 12'heff, 12'heee, 12'hdee, 12'hddd, 12'hccd, 12'hbad, 12'ha9c, 12'h98c, 12'h88b, 12'h98c, 12'ha9c, 12'hbad, 12'hbbd, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hdce, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'heee, 12'hfef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hedd, 12'hccb, 12'h999, 12'h777, 12'h655, 12'h555, 12'h544, 12'h434, 12'h444, 12'h545, 12'h545, 12'h445, 12'h446, 12'h556, 12'h557, 12'h789, 12'h99b, 12'hbbc, 12'hbbd, 12'hccd, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcce, 12'hccd, 12'hccd, 12'hbbc, 12'haac, 12'h9ab, 12'h99a, 12'h89a, 12'h99a, 12'h99a, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h66a, 
12'h669, 12'h559, 12'h448, 12'h338, 12'h438, 12'h549, 12'h659, 12'h66a, 12'h88b, 12'haac, 12'hcbd, 12'hcce, 12'hddf, 12'heef, 12'heef, 12'heef, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heef, 12'heef, 12'heff, 12'heef, 12'heee, 12'hdee, 12'hdde, 12'hcce, 12'hbbe, 12'hbad, 12'ha9d, 12'ha9c, 12'ha8c, 12'ha9c, 12'hbad, 12'hbad, 12'hbbd, 12'hcbd, 12'hcbd, 12'hbbd, 12'hcbd, 12'hccd, 12'hdce, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hede, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'hfee, 12'heed, 12'hdcc, 12'hbaa, 12'h988, 12'h766, 12'h655, 12'h544, 12'h434, 12'h434, 12'h545, 12'h545, 12'h445, 12'h445, 12'h546, 12'h557, 12'h779, 12'h99a, 12'haac, 12'hbbc, 12'hccd, 12'hcde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcde, 12'hcde, 12'hcce, 12'hccd, 12'hbbd, 12'habc, 12'h9ab, 12'h99a, 12'h89a, 12'h99a, 12'h89a, 12'h89b, 12'h88b, 12'h88b, 12'h88b, 12'h78b, 12'h77b, 12'h77a, 12'h77b, 12'h77a, 
12'h77a, 12'h76a, 12'h66a, 12'h659, 12'h659, 12'h659, 12'h659, 12'h66a, 12'h77a, 12'h99c, 12'hbbd, 12'hcce, 12'hdce, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heee, 12'hdee, 12'hdde, 12'hcdd, 12'hccd, 12'hbbd, 12'hbad, 12'hbad, 12'hbad, 12'hbad, 12'hbad, 12'hbad, 12'hbbd, 12'hcbd, 12'hcbd, 12'hcbd, 12'hccd, 12'hcce, 12'hdce, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 
12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hddd, 12'hcbb, 12'haaa, 12'h877, 12'h655, 12'h545, 12'h544, 12'h544, 12'h434, 12'h434, 12'h434, 12'h435, 12'h446, 12'h557, 12'h778, 12'h88a, 12'haab, 12'hbbc, 12'hccd, 12'hcde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcde, 12'hcde, 12'hcce, 12'hccd, 12'hbcd, 12'habc, 12'haab, 12'h99b, 12'h89a, 12'h89a, 12'h89a, 12'h88b, 12'h88b, 12'h88b, 12'h77b, 12'h77b, 12'h77a, 12'h77b, 12'h88b, 12'h88b, 
12'h88b, 12'h88b, 12'h88b, 12'h88b, 12'h87b, 12'h77a, 12'h66a, 12'h659, 12'h66a, 12'h88b, 12'haad, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcdd, 12'hccd, 12'hcbd, 12'hbbe, 12'hbae, 12'hbbe, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcbd, 12'hcbd, 12'hcbd, 12'hcce, 12'hcce, 12'hdce, 12'hdde, 12'hddf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 
12'heee, 12'hfef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hedd, 12'hdcc, 12'hbbb, 12'h888, 12'h655, 12'h655, 12'h655, 12'h545, 12'h434, 12'h324, 12'h324, 12'h435, 12'h446, 12'h557, 12'h668, 12'h789, 12'h99b, 12'hbbc, 12'hccd, 12'hcce, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hcde, 12'hcde, 12'hcce, 12'hccd, 12'hbcd, 12'hbbc, 12'haab, 12'h99b, 12'h89a, 12'h88a, 12'h88a, 12'h88a, 12'h78b, 12'h77b, 12'h77a, 12'h77a, 12'h77a, 12'h77b, 12'h88b, 12'h88b, 
12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h88b, 12'h87b, 12'h76a, 12'h77a, 12'h88b, 12'ha9c, 12'haad, 12'hbbd, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hcbd, 12'hcbe, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcbe, 12'hcbe, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 
12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hedd, 12'hccc, 12'ha99, 12'h766, 12'h766, 12'h655, 12'h545, 12'h434, 12'h434, 12'h324, 12'h334, 12'h445, 12'h556, 12'h557, 12'h778, 12'h99a, 12'haac, 12'hbbd, 12'hccd, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hccd, 12'hbcd, 12'hbbc, 12'haab, 12'h99b, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h77a, 12'h77b, 12'h77b, 12'h77a, 12'h77a, 12'h77a, 12'h77b, 12'h77b, 
12'h88b, 12'h88c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h98c, 12'h98c, 12'h98c, 12'h99c, 12'ha9c, 12'haad, 12'hbad, 12'haad, 12'haad, 12'haad, 12'haac, 12'haac, 12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbe, 12'hcce, 12'hdce, 12'hdcf, 12'hdcf, 12'hdcf, 12'hdcf, 12'hdce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 
12'hfef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'heee, 12'hddd, 12'hbba, 12'h988, 12'h877, 12'h656, 12'h545, 12'h544, 12'h434, 12'h324, 12'h324, 12'h445, 12'h546, 12'h557, 12'h668, 12'h88a, 12'haab, 12'hbbc, 12'hccd, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hbcd, 12'hbbc, 12'haac, 12'h99b, 12'h89a, 12'h789, 12'h779, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77a, 12'h77b, 12'h77b, 
12'h87b, 12'h88c, 12'h98c, 12'h99c, 12'h99d, 12'ha9d, 12'ha9d, 12'ha9d, 12'ha9d, 12'h99c, 12'h99c, 12'ha9d, 12'haad, 12'haad, 12'haad, 12'haad, 12'ha9c, 12'ha9c, 12'ha9c, 12'haad, 12'haad, 12'hbad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcbe, 12'hcce, 12'hcce, 12'hdce, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hddf, 12'hdce, 12'hdce, 12'hdce, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heef, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'hfee, 12'hedd, 12'hccc, 12'haa9, 12'h988, 12'h766, 12'h555, 12'h545, 12'h545, 12'h434, 12'h334, 12'h435, 12'h446, 12'h556, 12'h667, 12'h779, 12'h99b, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hcde, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hbcd, 12'hbbd, 12'haac, 12'h9ab, 12'h89a, 12'h779, 12'h669, 12'h669, 12'h669, 12'h66a, 12'h66a, 12'h77a, 12'h77a, 12'h77b, 12'h77b, 12'h77b, 
12'h77b, 12'h88b, 12'h88c, 12'h98c, 12'h99c, 12'ha9d, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbae, 12'hbae, 12'hbad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbad, 12'hbbd, 12'hbbe, 12'hcbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hedf, 12'hedf, 12'hedf, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hddc, 12'hcbb, 12'ha99, 12'h776, 12'h655, 12'h655, 12'h555, 12'h444, 12'h434, 12'h445, 12'h446, 12'h546, 12'h557, 12'h778, 12'h88a, 12'haab, 12'hbbc, 12'hbcd, 12'hccd, 12'hcce, 12'hcde, 12'hcde, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbbd, 12'haac, 12'h9ab, 12'h89a, 12'h679, 12'h568, 12'h558, 12'h459, 12'h559, 12'h569, 12'h66a, 12'h77a, 12'h77b, 12'h77b, 12'h77b, 
12'h87b, 12'h88b, 12'h88c, 12'h88c, 12'h99c, 12'h99d, 12'ha9d, 12'haad, 12'haad, 12'haae, 12'hbae, 12'hbae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbae, 12'hbae, 12'hbad, 12'hbad, 12'hbad, 12'hbae, 12'hbbe, 12'hcbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'hfef, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hedd, 12'hdcc, 12'hbaa, 12'h988, 12'h766, 12'h666, 12'h655, 12'h545, 12'h445, 12'h545, 12'h446, 12'h546, 12'h556, 12'h668, 12'h889, 12'h99a, 12'haac, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbbd, 12'habc, 12'h9ab, 12'h89a, 12'h779, 12'h568, 12'h458, 12'h448, 12'h458, 12'h559, 12'h569, 12'h66a, 12'h77a, 12'h77b, 12'h88b, 
12'h88b, 12'h88c, 12'h88c, 12'h88c, 12'h98c, 12'h99c, 12'h99d, 12'ha9d, 12'ha9d, 12'haad, 12'haae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbad, 12'hbae, 12'hbae, 12'hbbe, 12'hcbe, 12'hccf, 12'hddf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'hdde, 12'hdde, 12'hdde, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hedd, 12'hccc, 12'haa9, 12'h887, 12'h766, 12'h655, 12'h655, 12'h555, 12'h545, 12'h545, 12'h445, 12'h546, 12'h667, 12'h778, 12'h88a, 12'haab, 12'hbbc, 12'hbbd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'habc, 12'h9ac, 12'h89b, 12'h779, 12'h568, 12'h458, 12'h348, 12'h348, 12'h458, 12'h559, 12'h569, 12'h67a, 12'h77b, 12'h88b, 
12'h88b, 12'h99c, 12'h98c, 12'h88c, 12'h98c, 12'h98c, 12'h98c, 12'h98c, 12'h99d, 12'ha9d, 12'haad, 12'haae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'haae, 12'haae, 12'hbae, 12'hbae, 12'hbbe, 12'hccf, 12'hdcf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hdde, 12'hdde, 12'hede, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heee, 12'hddd, 12'hcbb, 12'ha99, 12'h877, 12'h766, 12'h666, 12'h666, 12'h556, 12'h555, 12'h445, 12'h446, 12'h557, 12'h668, 12'h889, 12'h99b, 12'haac, 12'hbbc, 12'hbbd, 12'hccd, 12'hccd, 12'hccd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habc, 12'haac, 12'h99b, 12'h78a, 12'h569, 12'h569, 12'h458, 12'h358, 12'h358, 12'h458, 12'h559, 12'h669, 12'h77a, 12'h88b, 
12'h88b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99d, 12'ha9d, 12'haad, 12'haad, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbae, 12'hbbe, 12'hbbe, 12'hccf, 12'hdcf, 12'hddf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'hedf, 12'hedf, 12'hedf, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'heed, 12'hddc, 12'hbbb, 12'h988, 12'h877, 12'h777, 12'h767, 12'h666, 12'h556, 12'h545, 12'h445, 12'h546, 12'h667, 12'h779, 12'h99a, 12'haab, 12'haac, 12'hbbc, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'haac, 12'h99b, 12'h88a, 12'h679, 12'h679, 12'h568, 12'h458, 12'h458, 12'h458, 12'h458, 12'h569, 12'h67a, 12'h77a, 
12'h88b, 12'h89b, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'h99c, 12'ha9d, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbae, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hccf, 12'hdcf, 12'hddf, 12'hddf, 12'hddf, 12'hede, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heed, 12'hdcc, 12'haaa, 12'h988, 12'h888, 12'h878, 12'h777, 12'h666, 12'h556, 12'h445, 12'h446, 12'h557, 12'h778, 12'h889, 12'h99a, 12'h99b, 12'haac, 12'hbbc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'hbbd, 12'hbbd, 12'habd, 12'habc, 12'h9ac, 12'h89b, 12'h78a, 12'h679, 12'h569, 12'h468, 12'h458, 12'h458, 12'h458, 12'h568, 12'h679, 12'h77a, 
12'h88b, 12'h89b, 12'h99b, 12'h99c, 12'h99c, 12'h9ac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hfee, 12'hedd, 12'hccb, 12'hbaa, 12'ha99, 12'h988, 12'h888, 12'h777, 12'h666, 12'h556, 12'h556, 12'h557, 12'h668, 12'h778, 12'h889, 12'h89a, 12'h99b, 12'haac, 12'habc, 12'habc, 12'hbbd, 12'habc, 12'habc, 12'habc, 12'habd, 12'habd, 12'habd, 12'habd, 12'haac, 12'h99b, 12'h78a, 12'h679, 12'h568, 12'h468, 12'h458, 12'h458, 12'h468, 12'h569, 12'h679, 12'h78a, 
12'h89b, 12'h99b, 12'h99c, 12'h9ac, 12'haac, 12'haac, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hbbe, 12'hbbe, 12'hcbe, 12'hcce, 12'hcce, 12'hccf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hbbb, 12'ha99, 12'h989, 12'h888, 12'h777, 12'h667, 12'h656, 12'h557, 12'h657, 12'h668, 12'h778, 12'h779, 12'h88a, 12'h99b, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'haac, 12'habd, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h89b, 12'h789, 12'h578, 12'h468, 12'h468, 12'h568, 12'h568, 12'h578, 12'h679, 12'h78a, 
12'h89a, 12'h99b, 12'h9ab, 12'haac, 12'haac, 12'haac, 12'habd, 12'habd, 12'habd, 12'haad, 12'haad, 12'haad, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbe, 12'hbbe, 12'hbbe, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hccc, 12'hbba, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h767, 12'h667, 12'h557, 12'h557, 12'h667, 12'h678, 12'h779, 12'h88a, 12'h99b, 12'haab, 12'haac, 12'haac, 12'h9ac, 12'h9ac, 12'haac, 12'habc, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h89b, 12'h78a, 12'h679, 12'h678, 12'h578, 12'h578, 12'h568, 12'h578, 12'h679, 12'h679, 
12'h78a, 12'h89b, 12'h9ab, 12'haac, 12'habc, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hddf, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'hddd, 12'hcbb, 12'hbaa, 12'haaa, 12'h999, 12'h989, 12'h888, 12'h667, 12'h556, 12'h556, 12'h557, 12'h567, 12'h678, 12'h88a, 12'h99b, 12'h99b, 12'h9ab, 12'h9ac, 12'h9ab, 12'h9ab, 12'h9ac, 12'haac, 12'habc, 12'habd, 12'habc, 12'h9ac, 12'h99b, 12'h89a, 12'h789, 12'h689, 12'h679, 12'h678, 12'h578, 12'h568, 12'h578, 12'h679, 
12'h789, 12'h89a, 12'h9ab, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'heee, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddc, 12'hccc, 12'hbbb, 12'haaa, 12'ha9a, 12'h999, 12'h878, 12'h667, 12'h557, 12'h557, 12'h557, 12'h668, 12'h779, 12'h88a, 12'h99a, 12'h99b, 12'h99b, 12'h99b, 12'h99b, 12'h9ab, 12'haac, 12'haac, 12'habd, 12'habd, 12'haac, 12'h9ac, 12'h99b, 12'h89a, 12'h789, 12'h789, 12'h679, 12'h679, 12'h678, 12'h679, 12'h679, 
12'h78a, 12'h89a, 12'h99b, 12'h9ac, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'hdee, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hbbb, 12'hbab, 12'haaa, 12'h999, 12'h888, 12'h778, 12'h667, 12'h668, 12'h668, 12'h779, 12'h889, 12'h88a, 12'h88a, 12'h89a, 12'h89b, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'habc, 12'habc, 12'habd, 12'habc, 12'h9ac, 12'h89b, 12'h89a, 12'h78a, 12'h78a, 12'h789, 12'h679, 12'h679, 12'h789, 
12'h78a, 12'h89a, 12'h89b, 12'h9ab, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heed, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'h99a, 12'h889, 12'h778, 12'h778, 12'h778, 12'h779, 12'h779, 12'h789, 12'h88a, 12'h88a, 12'h88a, 12'h89a, 12'h99b, 12'h9ab, 12'haac, 12'haac, 12'habc, 12'habd, 12'hbbd, 12'haac, 12'h9ab, 12'h99b, 12'h89b, 12'h89a, 12'h88a, 12'h78a, 12'h78a, 12'h78a, 
12'h78a, 12'h89a, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heee, 12'heee, 12'hddd, 12'hdcc, 12'hccc, 12'hbbb, 12'haab, 12'h99a, 12'h999, 12'h889, 12'h889, 12'h779, 12'h779, 12'h779, 12'h789, 12'h789, 12'h88a, 12'h88a, 12'h89b, 12'h99b, 12'h9ac, 12'haac, 12'habc, 12'habd, 12'hbbd, 12'habc, 12'habc, 12'haac, 12'h9ac, 12'h9ab, 12'h99b, 12'h89b, 12'h89b, 12'h89b, 
12'h89b, 12'h89b, 12'h99b, 12'h99b, 12'h9ac, 12'haac, 12'haac, 12'habc, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcde, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddf, 12'hddf, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'haaa, 12'haaa, 12'h99a, 12'h889, 12'h889, 12'h789, 12'h789, 12'h789, 12'h889, 12'h88a, 12'h89a, 12'h99b, 12'h9ab, 12'haac, 12'habc, 12'hbbc, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'haac, 12'haac, 12'h9ac, 12'h99b, 12'h99b, 12'h99b, 
12'h99b, 12'h99b, 12'h9ac, 12'h9ac, 12'haac, 12'haac, 12'habc, 12'habc, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcde, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hbbc, 12'hbbb, 12'haab, 12'h99a, 12'h99a, 12'h889, 12'h889, 12'h889, 12'h889, 12'h88a, 12'h89a, 12'h99b, 12'h9ab, 12'haac, 12'habc, 12'hbbd, 12'hbcd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'haac, 12'haac, 12'haac, 12'haac, 
12'haac, 12'haac, 12'haac, 12'haac, 12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'heee, 12'hdee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdef, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hede, 12'hddd, 12'hdcd, 12'hccc, 12'hbbc, 12'hbbb, 12'haab, 12'haaa, 12'h99a, 12'h99a, 12'h89a, 12'h89a, 12'h99a, 12'h99a, 12'h9ab, 12'haac, 12'hbbc, 12'hbcd, 12'hccd, 12'hccd, 12'hbce, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'habd, 12'habd, 12'habd, 
12'habd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hccd, 12'hbcd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbcd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hede, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heee, 12'heef, 12'heef, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hbbc, 12'hbbb, 12'haab, 12'haab, 12'haaa, 12'h9aa, 12'h99a, 12'h9ab, 12'haab, 12'habc, 12'hbbc, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hbbe, 12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 
12'hbbd, 12'hbbd, 12'hbbd, 12'hbbd, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heee, 12'heef, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hccc, 12'hbbc, 12'hbbb, 12'habb, 12'haab, 12'haab, 12'habb, 12'hbbc, 12'hbcc, 12'hccd, 12'hcde, 12'hcde, 12'hcde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hcdd, 12'hccc, 12'hccc, 12'hbbc, 12'hbbc, 12'hbbc, 12'hbcc, 12'hccd, 12'hccd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hcce, 12'hcce, 12'hcce, 12'hcce, 
12'hcce, 12'hcce, 12'hcce, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hccd, 12'hccc, 12'hccc, 12'hccd, 12'hccd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heef, 12'heef, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'heff, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 
12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 
12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hdde, 12'hdde, 
12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hcdd, 12'hddd, 12'hddd, 12'hcdd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'hdde, 12'hdde, 12'hdee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'heef, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 
12'heee, 12'heee, 12'heee, 12'hdee, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccd, 12'hccd, 12'hccd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hccd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 
12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hdde, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hdde, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h999, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h444, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h888, 12'h555, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h444, 12'h000, 12'h000, 12'h000, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h000, 12'h000, 12'h333, 12'h777, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h999, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h555, 12'h333, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'hdec, 12'hdec, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h7a2, 12'h6a0, 12'h6a0, 12'h8a4, 12'hddc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'hcdb, 12'hcdb, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h7a0, 12'h6a0, 12'h6a0, 12'h7a3, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hcda, 12'h9b7, 12'h9b7, 12'hbc9, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h8a4, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h7a2, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h000, 12'h555, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h000, 12'h444, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'hbca, 12'hbca, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'hded, 12'hfff, 12'hfff, 12'hbbb, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'h999, 12'h000, 12'h000, 12'h000, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h9b6, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'hfff, 12'h333, 12'h000, 12'h000, 12'h000, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'h777, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'h444, 12'h000, 12'h000, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hddd, 12'h555, 12'h000, 12'h333, 12'h999, 12'hfff, 12'hfff, 12'haaa, 12'h111, 12'h000, 12'h666, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h8a4, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'hcdc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbca, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9c7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a3, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbca, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hab7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h444, 12'h555, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbca, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h666, 12'h555, 12'h777, 12'hddd, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h555, 12'h000, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h000, 12'h000, 12'h000, 12'h000, 12'h666, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbca, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'h9b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'h000, 12'h000, 12'h444, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h777, 12'h999, 12'heee, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'hbca, 12'hac8, 12'hac9, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hded, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h9b6, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'hac8, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h9b6, 12'h8b5, 12'hac9, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hbca, 12'h8b5, 12'h7a0, 12'h6a0, 12'h7a1, 12'h9b6, 12'hcdb, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a3, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'h8b5, 12'hefe, 12'hfff, 12'hfff, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h6a0, 12'h7a0, 12'h6a0, 12'h7a3, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hded, 12'hded, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h9b6, 12'h6a0, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a0, 12'h7a0, 12'h6a0, 12'hbc9, 12'hfff, 12'hded, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'h8a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h8b5, 12'h7a0, 12'h6a0, 12'h6a0, 12'h7a1, 12'h9b6, 12'hefe, 12'hfff, 12'hfff, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'hac8, 12'hac9, 12'hded, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hefe, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'hbc9, 12'hbc9, 12'hdec, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h9b7, 12'h6a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a0, 12'h6a0, 12'h8b6, 12'hbda, 12'hac7, 12'h8a3, 12'h9b7, 12'hbc9, 12'hcdb, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h9b6, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'hbda, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hffe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'hac8, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h8a4, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'h7a0, 12'h7a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h8b5, 12'hcda, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hdec, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a3, 12'hffe, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hbda, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h6a0, 12'h6a0, 12'hbca, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbca, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbca, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hac8, 12'h6a0, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'h9b7, 12'heed, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'hbc9, 12'hac8, 12'hac8, 12'hbda, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hac9, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'hac8, 12'h6a0, 12'h8a3, 12'h7a2, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a3, 12'h7a3, 12'h9b6, 12'hdec, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'hefe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 
12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h8b5, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h7a3, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hbc9, 12'hac7, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'h9b7, 12'h6a0, 12'h8b4, 12'h7a3, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'h8b5, 12'h8b5, 12'hdec, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hac7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 
12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9c7, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hac8, 12'hac8, 12'hac7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a3, 12'h7a0, 12'h8b5, 12'hdec, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 
12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h8a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'hded, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h8b5, 12'h7a2, 12'hac8, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hefe, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h8b4, 12'hddc, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'heee, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 
12'h7a1, 12'hefe, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'hbda, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbca, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hac8, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hded, 12'h8a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hddc, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hded, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hdec, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hac8, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hbc9, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hcdc, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'hac9, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hffe, 12'hfff, 12'hfff, 12'hdec, 12'h8b4, 12'h6a0, 12'h7a0, 12'h7a2, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hddc, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'hcdb, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbca, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'hcdb, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hded, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hbda, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'heee, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h7a1, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hefe, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h9b6, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h8b4, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hffe, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hac8, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hac8, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hffe, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hac8, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'heed, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hbc9, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hcdb, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a3, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'hefe, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hac7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hbc9, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'hefe, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'h8b4, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hefe, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hddd, 12'h222, 12'h000, 12'h333, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h9b6, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hefe, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'h888, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'hbbb, 12'h000, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'heee, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbca, 12'hfff, 12'hfff, 12'hfff, 12'h111, 12'h000, 12'h000, 12'hccc, 12'hfff, 12'hddd, 12'h333, 12'h000, 12'h444, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'heed, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdc, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'h333, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a3, 12'hded, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hcdb, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hefe, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 12'hfff, 12'hfff, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbca, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbca, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 
12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hefe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 
12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b5, 12'hac7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hded, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'heee, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'h444, 12'h000, 12'h000, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'h999, 12'h666, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 
12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a3, 12'hac8, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hded, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdc, 12'hfff, 12'hfff, 12'hfff, 12'h555, 12'h000, 12'h000, 12'hddd, 12'hfff, 12'hfff, 12'hddd, 12'h000, 12'h000, 12'h888, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 
12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'hbc9, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hded, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h000, 12'h000, 12'h666, 12'heee, 12'heee, 12'h888, 12'h000, 12'h000, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 
12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'hac9, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'h666, 12'h000, 12'h000, 12'h000, 12'h222, 12'h000, 12'h000, 12'h222, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 
12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbca, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b5, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h999, 12'h777, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hcdc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hac7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h8a4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hbda, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h9b7, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hddc, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbda, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hddc, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a0, 12'h7a3, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h8b5, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hdec, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a0, 12'h7a0, 12'hded, 12'hcdb, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'h9b5, 12'h7a0, 12'h7a2, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'h8a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hded, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h8b5, 12'h8b4, 12'h7a0, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h6a0, 12'h8b4, 12'hac9, 12'hdec, 12'hffe, 12'hfff, 12'heee, 12'hdec, 12'hbca, 12'h9b7, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hdec, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a0, 12'h8b4, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'h9b6, 12'h7a0, 12'h7a3, 12'h7a2, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hffe, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h8b5, 12'hac8, 12'h8b4, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'heed, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'h6a0, 12'h7a3, 12'h8a4, 12'h7a1, 12'h6a0, 12'h6a0, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'heee, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'hded, 12'hfff, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hac7, 12'h7a1, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcda, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hded, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a2, 12'h8b4, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b5, 12'hfff, 12'hfff, 12'heed, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hfff, 12'hfff, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbc9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b7, 12'hcda, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b6, 12'hfff, 12'heed, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'h8b5, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hefe, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'h9b6, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a3, 12'hfff, 12'hfff, 12'h9b6, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h6a0, 12'hcda, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b5, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b6, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a1, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hddc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'heed, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hbc9, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hffe, 12'hfff, 12'hbc9, 12'h7a3, 12'h8b3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 
12'h7a1, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbda, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a0, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac9, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h8b5, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac9, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcda, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a1, 12'heee, 12'hfff, 12'h8b5, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h7a3, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'heed, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 
12'h9b6, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8a4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h8b5, 12'h6a0, 12'h6a0, 12'h6a0, 12'h8b5, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h9b7, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h7a2, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'h9b7, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h8b5, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h7a1, 12'hcdb, 12'hfff, 12'hfff, 12'heed, 12'h8a4, 12'h6a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h8b4, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a0, 12'h6a0, 12'h7a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'h9b6, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 
12'hac7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h7a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hac7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hddc, 12'hcdb, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddc, 12'h7a4, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'h8a4, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'h7a2, 12'h7a0, 12'h7a1, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hac8, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'hac8, 12'hac8, 12'hbca, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'hbc9, 12'h7a3, 12'h7a1, 12'h7a0, 12'h8b4, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdb, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h8b4, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h8b5, 12'h7a0, 12'h7a0, 12'h9b6, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcdc, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 
12'hbca, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'hac8, 12'h7a1, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'h7a0, 12'hac8, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'h7a4, 12'h6a0, 12'h7a1, 
12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'hbca, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h6a0, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h6a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h6a0, 12'h7a2, 
12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac7, 12'h6a0, 12'h6a0, 12'h6a0, 12'h7a3, 12'hcdb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbca, 12'h8a4, 12'h6a0, 12'h6a0, 12'h6a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h8a4, 12'hac9, 12'heed, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'h9b7, 12'h6a0, 
12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h6a0, 12'h9b6, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hac8, 12'h6a0, 12'h7a0, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a1, 12'h7a0, 12'h6a0, 12'h9b7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h9b7, 12'h7a1, 12'h7a1, 12'h8a4, 12'h9b7, 12'heed, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 12'hcdb, 12'hcdc, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdec, 12'hbca, 12'h9b7, 12'h8b5, 12'h8b4, 12'h7a3, 12'h8a3, 12'h8b5, 12'hac8, 12'hbda, 12'hdec, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heed, 
12'hbda, 12'hac9, 12'hac8, 12'hac8, 12'hbda, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbca, 12'h8a3, 12'h6a0, 12'h7a0, 12'h7a0, 12'h7a0, 12'h6a0, 12'h6a0, 12'hac8, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hefe, 12'hefe, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hffe, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hbca, 12'h9b6, 12'h8b5, 12'h9b5, 12'hac9, 12'hded, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'heee, 12'hfff, 12'hddd, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'heee, 
12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hddd, 12'hccc, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hccc, 12'heee, 12'hccc, 12'hbbb, 12'hccc, 12'hddd, 12'heee, 12'hddd, 12'hbbb, 12'heee, 12'heee, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hccc, 12'heee, 12'hccc, 12'haaa, 12'hccc, 12'hbbb, 12'haaa, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'heee, 12'hccc, 12'hccc, 12'hddd, 12'hfff, 12'heee, 12'hccc, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hccc, 12'hddd, 12'heee, 12'heee, 12'hccc, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hddd, 12'hbbb, 12'hccc, 12'heee, 12'heee, 12'hccc, 12'heee, 12'hbbb, 12'haaa, 12'hddd, 12'hddd, 12'hddd, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hccc, 12'hfff, 12'hddd, 12'hccc, 12'heee, 12'hddd, 12'hfff, 12'hbbb, 12'heee, 12'hddd, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'heee, 12'heee, 12'hddd, 12'heee, 12'hfff, 12'heee, 12'hccc, 12'hddd, 12'hfff, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'hbbb, 12'hccc, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hddd, 12'heee, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hfff, 12'hddd, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'haaa, 12'hbbb, 12'heee, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hddd, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hfff, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'haaa, 12'hccc, 12'hddd, 12'hccc, 12'hccc, 12'hddd, 12'hccc, 12'haaa, 12'haaa, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hbbb, 12'h999, 12'hbbb, 12'hddd, 
12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hccc, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff};


	reg [11:0] pix_value; // the output pixel value according to the position and mode of the input
	reg [9:0]x_loc, y_loc; // x and y values
	reg [16:0]pix_val; // index of the pixel needed for the the output
	reg [11:0] D_in; // temporary reg
	always @(*)begin
		if (mode == 4'b1010)
			D_in<=12'hfff;
		else if (mode == 13)begin
			pix_val <= x + y * 640;
			D_in <= data[{pix_val}];
		end else begin
		pix_val <= 6400 * mode +((x%80) + ((y%80) * 80));
		D_in <= data[{pix_val}];
	end
//	else begin
//		if (mode==11) begin
//				pix_val <= 6400*2 * (mode%10-1) +((x%160) + ((y%80) * 80));
//				D_in <= background[{pix_val}];
//		end
//		else begin
//				pix_val <= 6400*2 * (mode%10-1) +((x%160) + ((y%80) * 80));
//				D_in <= background[{pix_val}];
//		end
//end
	end
	assign out = D_in;

endmodule
