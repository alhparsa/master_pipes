`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:50:28 01/03/2019 
// Design Name: 
// Module Name:    pipesmod 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pipesmod(input [9:0] x,
                input[9:0] y,
                output [7:0] D_in
					 //output [9:0] x_o,
					 //output {9:0] y_o
                );
	 
	
 //wire [9:0] x_loc = 160 + 80 * (x % 3);
 //wire [9:0] y_loc = 80 + 80 * (y / 3);
 wire [9:0] x_loc = (x-200) % 80;
 wire [9:0] y_loc = (y-119) %80;
	 
	 //assign x_o = x;
	 //assign y_o = y;
	
	 wire [9:0] elementnum = y_loc*80 + x_loc;
	
	parameter data = {8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe
,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe
,8'hfe,8'hfe,8'hfd,8'hfd,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbd,8'hfd,8'hfe,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hbd,8'hbd,8'hbd,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc
,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc
,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc
,8'hbc,8'hbc,8'hbc,8'hbc,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb
,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'h7b,8'h7a,8'h7a
,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h30,8'hbb,8'hbc,8'hfd,8'hfe,8'hff,8'hff,8'hff
,8'h79,8'h79,8'h79,8'h79,8'h78,8'h38,8'h38,8'h38,8'h38,8'h38,8'h78,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h78,8'h78,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h39,8'h39,8'h39,8'h39,8'h39,8'h38
,8'h38,8'h38,8'h38,8'h78,8'h78,8'h79,8'hbc,8'hfe,8'hff,8'hff,8'h39,8'h39,8'h39,8'h38
,8'h38,8'h38,8'h38,8'h39,8'h38,8'h38,8'h79,8'h79,8'h38,8'h38,8'h79,8'h79,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h39,8'h39,8'h39,8'h39,8'h39,8'h3a
,8'h3a,8'h3a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h78,8'h38,8'h38,8'h38
,8'h38,8'h78,8'h78,8'h78,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h79
,8'h38,8'h38,8'h38,8'hbc,8'hfe,8'hff,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h39,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h7a,8'h7a,8'h79,8'h7a,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a
,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h39,8'h39,8'h39,8'h39,8'h79,8'h79,8'h79
,8'h78,8'h38,8'h38,8'h38,8'h38,8'h79,8'h79,8'h79,8'h31,8'h79,8'h38,8'h38,8'h38,8'h32
,8'hbc,8'hfd,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h38,8'h78,8'h78
,8'h38,8'h38,8'h38,8'h78,8'h79,8'h39,8'h39,8'h38,8'h38,8'h39,8'h39,8'h79,8'h39,8'h38
,8'h38,8'h38,8'h39,8'h39,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h39,8'h39,8'h39,8'h79,8'h79,8'h79,8'h79,8'h79,8'h38,8'h38,8'h38,8'h38
,8'h78,8'h78,8'h38,8'h38,8'h7a,8'h7a,8'h70,8'h39,8'h3a,8'h39,8'h7a,8'hbb,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h38,8'h38,8'h38,8'h39
,8'h39,8'h3a,8'h3a,8'h3a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h38,8'h78,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h7a
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h38,8'h78,8'h79,8'h78,8'h78,8'h78,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h39,8'h79
,8'h70,8'h78,8'h78,8'h38,8'h38,8'h78,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h39,8'h39,8'h70,8'h78,8'h39,8'h38
,8'h79,8'hbb,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h3a,8'h79,8'h78,8'h38,8'h38,8'h32,8'hbb,8'hbd,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h3a,8'h79,8'h78,8'h38,8'h79,8'hbb,8'hfd,8'hfe,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h3a,8'h79,8'h78,8'h78
,8'hbb,8'hbd,8'hfe,8'hff,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h78,8'h78,8'h78
,8'h78,8'h38,8'h38,8'h78,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h38,8'h78,8'h78,8'h78,8'h38,8'h38,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h7a,8'h7a,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h38,8'h38,8'h79,8'h79
,8'h79,8'h78,8'h78,8'h38,8'h78,8'h78,8'h38,8'h39,8'hb3,8'hbc,8'hfe,8'hff,8'hff,8'hff
,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79,8'h71,8'h71,8'h39,8'h39,8'h39,8'h39,8'h39,8'h39
,8'h39,8'h79,8'h39,8'h39,8'h38,8'h38,8'h38,8'h38,8'h39,8'h39,8'h39,8'h39,8'h39,8'h39
,8'h39,8'h39,8'h39,8'h39,8'h78,8'h78,8'h38,8'h38,8'h38,8'h78,8'h78,8'h78,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h79,8'h7a
,8'h7a,8'hbb,8'hbc,8'hbc,8'hfd,8'hfe,8'hff,8'hff,8'hff,8'hff,8'h39,8'h39,8'h79,8'h79
,8'h79,8'h7a,8'h7a,8'h79,8'h39,8'h7a,8'h7a,8'h7a,8'h3a,8'h39,8'h3a,8'h7a,8'h7a,8'h7a
,8'h7a,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h3a,8'h3a,8'h7a,8'h7a,8'h7a,8'h3a
,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a
,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'hba
,8'hbb,8'hbb,8'hbb,8'hbb,8'hbc,8'hbc,8'hbc,8'hbc,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbd,8'hbd,8'hbd
,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd
,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd
,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe
,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe
,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff};
	
 /*
    reg [6399:0] pixel_in [7:0] = {8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe
,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe
,8'hfe,8'hfe,8'hfd,8'hfd,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbd,8'hfd,8'hfe,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hbd,8'hbd,8'hbd,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc
,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc
,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc
,8'hbc,8'hbc,8'hbc,8'hbc,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb
,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'h7b,8'h7a,8'h7a
,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h30,8'hbb,8'hbc,8'hfd,8'hfe,8'hff,8'hff,8'hff
,8'h79,8'h79,8'h79,8'h79,8'h78,8'h38,8'h38,8'h38,8'h38,8'h38,8'h78,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h78,8'h78,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h39,8'h39,8'h39,8'h39,8'h39,8'h38
,8'h38,8'h38,8'h38,8'h78,8'h78,8'h79,8'hbc,8'hfe,8'hff,8'hff,8'h39,8'h39,8'h39,8'h38
,8'h38,8'h38,8'h38,8'h39,8'h38,8'h38,8'h79,8'h79,8'h38,8'h38,8'h79,8'h79,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h39,8'h39,8'h39,8'h39,8'h39,8'h3a
,8'h3a,8'h3a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h78,8'h38,8'h38,8'h38
,8'h38,8'h78,8'h78,8'h78,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h79
,8'h38,8'h38,8'h38,8'hbc,8'hfe,8'hff,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h39,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h7a,8'h7a,8'h79,8'h7a,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a
,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h39,8'h39,8'h39,8'h39,8'h79,8'h79,8'h79
,8'h78,8'h38,8'h38,8'h38,8'h38,8'h79,8'h79,8'h79,8'h31,8'h79,8'h38,8'h38,8'h38,8'h32
,8'hbc,8'hfd,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h38,8'h78,8'h78
,8'h38,8'h38,8'h38,8'h78,8'h79,8'h39,8'h39,8'h38,8'h38,8'h39,8'h39,8'h79,8'h39,8'h38
,8'h38,8'h38,8'h39,8'h39,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h39,8'h39,8'h39,8'h79,8'h79,8'h79,8'h79,8'h79,8'h38,8'h38,8'h38,8'h38
,8'h78,8'h78,8'h38,8'h38,8'h7a,8'h7a,8'h70,8'h39,8'h3a,8'h39,8'h7a,8'hbb,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h38,8'h38,8'h38,8'h39
,8'h39,8'h3a,8'h3a,8'h3a,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h38,8'h78,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h7a
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h38,8'h78,8'h79,8'h78,8'h78,8'h78,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h39,8'h79
,8'h70,8'h78,8'h78,8'h38,8'h38,8'h78,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h39,8'h39,8'h70,8'h78,8'h39,8'h38
,8'h79,8'hbb,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h3a,8'h79,8'h78,8'h38,8'h38,8'h32,8'hbb,8'hbd,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h3a,8'h79,8'h78,8'h38,8'h79,8'hbb,8'hfd,8'hfe,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h3a,8'h79,8'h78,8'h78
,8'hbb,8'hbd,8'hfe,8'hff,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h78,8'h78,8'h78
,8'h78,8'h38,8'h38,8'h78,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h38,8'h78,8'h78,8'h78,8'h38,8'h38,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h7a,8'h7a,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h79,8'h79
,8'h79,8'h79,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h79,8'h79,8'h79,8'h38,8'h38,8'h79,8'h79
,8'h79,8'h78,8'h78,8'h38,8'h78,8'h78,8'h38,8'h39,8'hb3,8'hbc,8'hfe,8'hff,8'hff,8'hff
,8'h78,8'h78,8'h79,8'h79,8'h79,8'h79,8'h71,8'h71,8'h39,8'h39,8'h39,8'h39,8'h39,8'h39
,8'h39,8'h79,8'h39,8'h39,8'h38,8'h38,8'h38,8'h38,8'h39,8'h39,8'h39,8'h39,8'h39,8'h39
,8'h39,8'h39,8'h39,8'h39,8'h78,8'h78,8'h38,8'h38,8'h38,8'h78,8'h78,8'h78,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38
,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h38,8'h79,8'h7a
,8'h7a,8'hbb,8'hbc,8'hbc,8'hfd,8'hfe,8'hff,8'hff,8'hff,8'hff,8'h39,8'h39,8'h79,8'h79
,8'h79,8'h7a,8'h7a,8'h79,8'h39,8'h7a,8'h7a,8'h7a,8'h3a,8'h39,8'h3a,8'h7a,8'h7a,8'h7a
,8'h7a,8'h79,8'h79,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h3a,8'h3a,8'h7a,8'h7a,8'h7a,8'h3a
,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a
,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'hba
,8'hbb,8'hbb,8'hbb,8'hbb,8'hbc,8'hbc,8'hbc,8'hbc,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hbc,8'hbc,8'hbc,8'hbc,8'hbc,8'hbd,8'hbd,8'hbd
,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd
,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd
,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe
,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe
,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff
,8'hff,8'hff}; 
   */
assign D_in = 8'b1111_1111;
//assign D_in = data[elementnum];
//assign D_in = pixel_in[elementnum];
    //x_loc is 8 bits, y_loc is 8 bits, we want d out
	 


endmodule
